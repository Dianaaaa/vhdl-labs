// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.11.0.396.4
// Netlist written on Thu Nov 19 19:56:36 2020
//
// Verilog Description of module cpu2system
//

module cpu2system (clk, reset, akku_o);   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(7[8:18])
    input clk;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(8[13:16])
    input reset;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(9[13:18])
    output [8:0]akku_o;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(8[13:16])
    wire mem_0__7__N_83 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_0__7__N_83 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_1__7__N_88 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_1__7__N_88 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_2__7__N_91 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_2__7__N_91 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_3__7__N_94 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_3__7__N_94 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_4__7__N_97 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_4__7__N_97 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_5__7__N_100 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_5__7__N_100 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_6__7__N_103 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_6__7__N_103 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_8__7__N_109 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_8__7__N_109 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_9__7__N_112 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_9__7__N_112 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_10__7__N_115 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_10__7__N_115 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_11__7__N_118 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_11__7__N_118 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_12__7__N_121 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_12__7__N_121 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_13__7__N_124 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_13__7__N_124 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_14__7__N_127 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_14__7__N_127 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_16__7__N_133 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_16__7__N_133 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_17__7__N_136 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_17__7__N_136 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_18__7__N_139 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_18__7__N_139 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_19__7__N_142 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_19__7__N_142 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_20__7__N_145 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_20__7__N_145 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_21__7__N_148 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_21__7__N_148 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_22__7__N_151 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_22__7__N_151 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_24__7__N_157 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_24__7__N_157 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_25__7__N_160 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_25__7__N_160 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_26__7__N_163 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_26__7__N_163 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_27__7__N_166 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_27__7__N_166 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_28__7__N_169 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_28__7__N_169 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_29__7__N_172 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_29__7__N_172 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_30__7__N_175 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_30__7__N_175 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_32__7__N_181 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_32__7__N_181 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_33__7__N_184 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_33__7__N_184 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_34__7__N_187 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_34__7__N_187 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_35__7__N_190 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_35__7__N_190 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_36__7__N_193 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_36__7__N_193 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_37__7__N_196 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_37__7__N_196 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_38__7__N_199 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_38__7__N_199 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_40__7__N_205 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_40__7__N_205 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_41__7__N_208 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_41__7__N_208 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_42__7__N_211 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_42__7__N_211 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_43__7__N_214 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_43__7__N_214 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_44__7__N_217 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_44__7__N_217 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_45__7__N_220 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_45__7__N_220 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_46__7__N_223 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_46__7__N_223 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_48__7__N_229 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_48__7__N_229 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_49__7__N_232 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_49__7__N_232 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_50__7__N_235 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_50__7__N_235 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_51__7__N_238 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_51__7__N_238 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_52__7__N_241 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_52__7__N_241 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_53__7__N_244 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_53__7__N_244 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_54__7__N_247 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_54__7__N_247 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_56__7__N_253 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_56__7__N_253 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_57__7__N_256 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_57__7__N_256 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_58__7__N_259 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_58__7__N_259 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_59__7__N_262 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_59__7__N_262 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_60__7__N_265 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_60__7__N_265 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_61__7__N_268 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_61__7__N_268 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_62__7__N_271 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_62__7__N_271 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire GND_net, reset_c, akku_o_c_8, akku_o_c_7, akku_o_c_6, akku_o_c_5, 
        akku_o_c_4, akku_o_c_3, akku_o_c_2, akku_o_c_1, akku_o_c_0;
    wire [7:0]data;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(37[13:17])
    wire [5:0]pc_5__N_30;
    
    wire n1272;
    wire [5:0]address;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(24[9:16])
    
    wire n1287, n1295, n1290, n1292, n1289, n1286, n684, n681, 
        data_7__N_79, n1283, n1891, n1890, n1261, n1293, n1284, 
        n1296, n1260, VCC_net;
    
    IB reset_pad (.I(reset), .O(reset_c));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(9[13:18])
    IB clk_pad (.I(clk), .O(clk_c));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(8[13:16])
    OB akku_o_pad_0 (.I(akku_o_c_0), .O(akku_o[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_1 (.I(akku_o_c_1), .O(akku_o[1]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_2 (.I(akku_o_c_2), .O(akku_o[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_3 (.I(akku_o_c_3), .O(akku_o[3]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_4 (.I(akku_o_c_4), .O(akku_o[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_5 (.I(akku_o_c_5), .O(akku_o[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_6 (.I(akku_o_c_6), .O(akku_o[6]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_7 (.I(akku_o_c_7), .O(akku_o[7]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_8 (.I(akku_o_c_8), .O(akku_o[8]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    GSR GSR_INST (.GSR(reset_c));
    \sram64kx8("sram64kx8.dat")(1,13)  RAM (.address({address}), .mem_62__7__N_271(mem_62__7__N_271), 
            .data({data}), .mem_61__7__N_268(mem_61__7__N_268), .n1290(n1290), 
            .n1289(n1289), .n1283(n1283), .n1284(n1284), .n1293(n1293), 
            .mem_60__7__N_265(mem_60__7__N_265), .mem_59__7__N_262(mem_59__7__N_262), 
            .mem_58__7__N_259(mem_58__7__N_259), .mem_57__7__N_256(mem_57__7__N_256), 
            .mem_56__7__N_253(mem_56__7__N_253), .mem_54__7__N_247(mem_54__7__N_247), 
            .mem_53__7__N_244(mem_53__7__N_244), .mem_52__7__N_241(mem_52__7__N_241), 
            .mem_51__7__N_238(mem_51__7__N_238), .mem_50__7__N_235(mem_50__7__N_235), 
            .mem_49__7__N_232(mem_49__7__N_232), .mem_48__7__N_229(mem_48__7__N_229), 
            .mem_46__7__N_223(mem_46__7__N_223), .mem_45__7__N_220(mem_45__7__N_220), 
            .mem_44__7__N_217(mem_44__7__N_217), .mem_43__7__N_214(mem_43__7__N_214), 
            .mem_42__7__N_211(mem_42__7__N_211), .mem_41__7__N_208(mem_41__7__N_208), 
            .mem_40__7__N_205(mem_40__7__N_205), .mem_38__7__N_199(mem_38__7__N_199), 
            .mem_37__7__N_196(mem_37__7__N_196), .mem_36__7__N_193(mem_36__7__N_193), 
            .mem_35__7__N_190(mem_35__7__N_190), .mem_34__7__N_187(mem_34__7__N_187), 
            .mem_33__7__N_184(mem_33__7__N_184), .mem_32__7__N_181(mem_32__7__N_181), 
            .mem_30__7__N_175(mem_30__7__N_175), .mem_29__7__N_172(mem_29__7__N_172), 
            .mem_28__7__N_169(mem_28__7__N_169), .mem_27__7__N_166(mem_27__7__N_166), 
            .mem_26__7__N_163(mem_26__7__N_163), .mem_25__7__N_160(mem_25__7__N_160), 
            .mem_24__7__N_157(mem_24__7__N_157), .mem_22__7__N_151(mem_22__7__N_151), 
            .mem_21__7__N_148(mem_21__7__N_148), .mem_20__7__N_145(mem_20__7__N_145), 
            .mem_19__7__N_142(mem_19__7__N_142), .mem_18__7__N_139(mem_18__7__N_139), 
            .mem_17__7__N_136(mem_17__7__N_136), .mem_16__7__N_133(mem_16__7__N_133), 
            .mem_14__7__N_127(mem_14__7__N_127), .mem_13__7__N_124(mem_13__7__N_124), 
            .mem_12__7__N_121(mem_12__7__N_121), .mem_11__7__N_118(mem_11__7__N_118), 
            .mem_10__7__N_115(mem_10__7__N_115), .mem_9__7__N_112(mem_9__7__N_112), 
            .mem_8__7__N_109(mem_8__7__N_109), .mem_6__7__N_103(mem_6__7__N_103), 
            .mem_5__7__N_100(mem_5__7__N_100), .mem_4__7__N_97(mem_4__7__N_97), 
            .mem_3__7__N_94(mem_3__7__N_94), .mem_2__7__N_91(mem_2__7__N_91), 
            .mem_1__7__N_88(mem_1__7__N_88), .mem_0__7__N_83(mem_0__7__N_83), 
            .n1292(n1292), .n1296(n1296), .akku_o_c_0(akku_o_c_0), .data_7__N_79(data_7__N_79), 
            .n1891(n1891), .n684(n684), .n1272(n1272), .n1890(n1890), 
            .n1260(n1260), .n1261(n1261), .n1295(n1295), .n681(n681), 
            .n1287(n1287), .n1286(n1286), .akku_o_c_1(akku_o_c_1), .akku_o_c_2(akku_o_c_2), 
            .akku_o_c_3(akku_o_c_3), .akku_o_c_4(akku_o_c_4), .akku_o_c_5(akku_o_c_5), 
            .akku_o_c_6(akku_o_c_6), .akku_o_c_7(akku_o_c_7), .\pc_5__N_30[0] (pc_5__N_30[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(44[10:19])
    VLO i1 (.Z(GND_net));
    TSALL TSALL_INST (.TSALL(GND_net));
    CPU8BIT2 CPU (.akku_o_c_0(akku_o_c_0), .clk_c(clk_c), .reset_c(reset_c), 
            .n1891(n1891), .n1296(n1296), .n1290(n1290), .mem_12__7__N_121(mem_12__7__N_121), 
            .data_7__N_79(data_7__N_79), .pc_5__N_30({Open_0, Open_1, 
            Open_2, Open_3, Open_4, pc_5__N_30[0]}), .n1287(n1287), 
            .n1289(n1289), .mem_6__7__N_103(mem_6__7__N_103), .n1286(n1286), 
            .n1272(n1272), .mem_58__7__N_259(mem_58__7__N_259), .GND_net(GND_net), 
            .data({data}), .akku_o_c_6(akku_o_c_6), .akku_o_c_7(akku_o_c_7), 
            .akku_o_c_4(akku_o_c_4), .akku_o_c_5(akku_o_c_5), .akku_o_c_2(akku_o_c_2), 
            .akku_o_c_3(akku_o_c_3), .akku_o_c_1(akku_o_c_1), .address({address}), 
            .n1890(n1890), .akku_o_c_8(akku_o_c_8), .n1293(n1293), .mem_59__7__N_262(mem_59__7__N_262), 
            .mem_60__7__N_265(mem_60__7__N_265), .n681(n681), .mem_61__7__N_268(mem_61__7__N_268), 
            .mem_62__7__N_271(mem_62__7__N_271), .n1295(n1295), .n1283(n1283), 
            .mem_48__7__N_229(mem_48__7__N_229), .n1292(n1292), .mem_49__7__N_232(mem_49__7__N_232), 
            .mem_50__7__N_235(mem_50__7__N_235), .mem_51__7__N_238(mem_51__7__N_238), 
            .mem_52__7__N_241(mem_52__7__N_241), .mem_53__7__N_244(mem_53__7__N_244), 
            .mem_54__7__N_247(mem_54__7__N_247), .n1260(n1260), .mem_40__7__N_205(mem_40__7__N_205), 
            .mem_41__7__N_208(mem_41__7__N_208), .mem_42__7__N_211(mem_42__7__N_211), 
            .mem_43__7__N_214(mem_43__7__N_214), .mem_44__7__N_217(mem_44__7__N_217), 
            .mem_45__7__N_220(mem_45__7__N_220), .mem_46__7__N_223(mem_46__7__N_223), 
            .n1284(n1284), .mem_32__7__N_181(mem_32__7__N_181), .mem_33__7__N_184(mem_33__7__N_184), 
            .mem_34__7__N_187(mem_34__7__N_187), .mem_35__7__N_190(mem_35__7__N_190), 
            .mem_36__7__N_193(mem_36__7__N_193), .mem_37__7__N_196(mem_37__7__N_196), 
            .mem_38__7__N_199(mem_38__7__N_199), .n684(n684), .mem_24__7__N_157(mem_24__7__N_157), 
            .mem_25__7__N_160(mem_25__7__N_160), .mem_26__7__N_163(mem_26__7__N_163), 
            .mem_27__7__N_166(mem_27__7__N_166), .mem_28__7__N_169(mem_28__7__N_169), 
            .mem_29__7__N_172(mem_29__7__N_172), .mem_30__7__N_175(mem_30__7__N_175), 
            .n1261(n1261), .mem_16__7__N_133(mem_16__7__N_133), .mem_17__7__N_136(mem_17__7__N_136), 
            .mem_18__7__N_139(mem_18__7__N_139), .mem_19__7__N_142(mem_19__7__N_142), 
            .mem_20__7__N_145(mem_20__7__N_145), .mem_21__7__N_148(mem_21__7__N_148), 
            .mem_22__7__N_151(mem_22__7__N_151), .mem_8__7__N_109(mem_8__7__N_109), 
            .mem_9__7__N_112(mem_9__7__N_112), .mem_10__7__N_115(mem_10__7__N_115), 
            .mem_5__7__N_100(mem_5__7__N_100), .mem_57__7__N_256(mem_57__7__N_256), 
            .mem_56__7__N_253(mem_56__7__N_253), .mem_4__7__N_97(mem_4__7__N_97), 
            .mem_3__7__N_94(mem_3__7__N_94), .mem_2__7__N_91(mem_2__7__N_91), 
            .mem_1__7__N_88(mem_1__7__N_88), .mem_0__7__N_83(mem_0__7__N_83), 
            .mem_14__7__N_127(mem_14__7__N_127), .mem_13__7__N_124(mem_13__7__N_124), 
            .mem_11__7__N_118(mem_11__7__N_118));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(43[10:18])
    VHI i2042 (.Z(VCC_net));
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module \sram64kx8("sram64kx8.dat")(1,13) 
//

module \sram64kx8("sram64kx8.dat")(1,13)  (address, mem_62__7__N_271, data, 
            mem_61__7__N_268, n1290, n1289, n1283, n1284, n1293, 
            mem_60__7__N_265, mem_59__7__N_262, mem_58__7__N_259, mem_57__7__N_256, 
            mem_56__7__N_253, mem_54__7__N_247, mem_53__7__N_244, mem_52__7__N_241, 
            mem_51__7__N_238, mem_50__7__N_235, mem_49__7__N_232, mem_48__7__N_229, 
            mem_46__7__N_223, mem_45__7__N_220, mem_44__7__N_217, mem_43__7__N_214, 
            mem_42__7__N_211, mem_41__7__N_208, mem_40__7__N_205, mem_38__7__N_199, 
            mem_37__7__N_196, mem_36__7__N_193, mem_35__7__N_190, mem_34__7__N_187, 
            mem_33__7__N_184, mem_32__7__N_181, mem_30__7__N_175, mem_29__7__N_172, 
            mem_28__7__N_169, mem_27__7__N_166, mem_26__7__N_163, mem_25__7__N_160, 
            mem_24__7__N_157, mem_22__7__N_151, mem_21__7__N_148, mem_20__7__N_145, 
            mem_19__7__N_142, mem_18__7__N_139, mem_17__7__N_136, mem_16__7__N_133, 
            mem_14__7__N_127, mem_13__7__N_124, mem_12__7__N_121, mem_11__7__N_118, 
            mem_10__7__N_115, mem_9__7__N_112, mem_8__7__N_109, mem_6__7__N_103, 
            mem_5__7__N_100, mem_4__7__N_97, mem_3__7__N_94, mem_2__7__N_91, 
            mem_1__7__N_88, mem_0__7__N_83, n1292, n1296, akku_o_c_0, 
            data_7__N_79, n1891, n684, n1272, n1890, n1260, n1261, 
            n1295, n681, n1287, n1286, akku_o_c_1, akku_o_c_2, akku_o_c_3, 
            akku_o_c_4, akku_o_c_5, akku_o_c_6, akku_o_c_7, \pc_5__N_30[0] );
    input [5:0]address;
    input mem_62__7__N_271;
    output [7:0]data;
    input mem_61__7__N_268;
    output n1290;
    output n1289;
    output n1283;
    output n1284;
    output n1293;
    input mem_60__7__N_265;
    input mem_59__7__N_262;
    input mem_58__7__N_259;
    input mem_57__7__N_256;
    input mem_56__7__N_253;
    input mem_54__7__N_247;
    input mem_53__7__N_244;
    input mem_52__7__N_241;
    input mem_51__7__N_238;
    input mem_50__7__N_235;
    input mem_49__7__N_232;
    input mem_48__7__N_229;
    input mem_46__7__N_223;
    input mem_45__7__N_220;
    input mem_44__7__N_217;
    input mem_43__7__N_214;
    input mem_42__7__N_211;
    input mem_41__7__N_208;
    input mem_40__7__N_205;
    input mem_38__7__N_199;
    input mem_37__7__N_196;
    input mem_36__7__N_193;
    input mem_35__7__N_190;
    input mem_34__7__N_187;
    input mem_33__7__N_184;
    input mem_32__7__N_181;
    input mem_30__7__N_175;
    input mem_29__7__N_172;
    input mem_28__7__N_169;
    input mem_27__7__N_166;
    input mem_26__7__N_163;
    input mem_25__7__N_160;
    input mem_24__7__N_157;
    input mem_22__7__N_151;
    input mem_21__7__N_148;
    input mem_20__7__N_145;
    input mem_19__7__N_142;
    input mem_18__7__N_139;
    input mem_17__7__N_136;
    input mem_16__7__N_133;
    input mem_14__7__N_127;
    input mem_13__7__N_124;
    input mem_12__7__N_121;
    input mem_11__7__N_118;
    input mem_10__7__N_115;
    input mem_9__7__N_112;
    input mem_8__7__N_109;
    input mem_6__7__N_103;
    input mem_5__7__N_100;
    input mem_4__7__N_97;
    input mem_3__7__N_94;
    input mem_2__7__N_91;
    input mem_1__7__N_88;
    input mem_0__7__N_83;
    output n1292;
    output n1296;
    input akku_o_c_0;
    input data_7__N_79;
    input n1891;
    output n684;
    output n1272;
    input n1890;
    output n1260;
    output n1261;
    output n1295;
    output n681;
    output n1287;
    output n1286;
    input akku_o_c_1;
    input akku_o_c_2;
    input akku_o_c_3;
    input akku_o_c_4;
    input akku_o_c_5;
    input akku_o_c_6;
    input akku_o_c_7;
    output \pc_5__N_30[0] ;
    
    wire mem_62__7__N_271 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_62__7__N_271 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_61__7__N_268 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_61__7__N_268 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_60__7__N_265 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_60__7__N_265 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_59__7__N_262 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_59__7__N_262 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_58__7__N_259 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_58__7__N_259 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_57__7__N_256 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_57__7__N_256 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_56__7__N_253 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_56__7__N_253 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_55__7__N_250 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_55__7__N_250 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_54__7__N_247 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_54__7__N_247 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_53__7__N_244 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_53__7__N_244 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_52__7__N_241 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_52__7__N_241 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_51__7__N_238 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_51__7__N_238 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_50__7__N_235 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_50__7__N_235 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_49__7__N_232 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_49__7__N_232 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_48__7__N_229 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_48__7__N_229 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_47__7__N_226 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_47__7__N_226 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_46__7__N_223 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_46__7__N_223 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_45__7__N_220 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_45__7__N_220 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_44__7__N_217 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_44__7__N_217 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_43__7__N_214 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_43__7__N_214 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_42__7__N_211 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_42__7__N_211 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_41__7__N_208 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_41__7__N_208 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_40__7__N_205 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_40__7__N_205 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_39__7__N_202 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_39__7__N_202 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_38__7__N_199 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_38__7__N_199 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_37__7__N_196 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_37__7__N_196 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_36__7__N_193 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_36__7__N_193 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_35__7__N_190 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_35__7__N_190 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_34__7__N_187 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_34__7__N_187 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_33__7__N_184 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_33__7__N_184 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_32__7__N_181 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_32__7__N_181 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_31__7__N_178 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_31__7__N_178 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_30__7__N_175 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_30__7__N_175 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_29__7__N_172 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_29__7__N_172 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_28__7__N_169 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_28__7__N_169 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_27__7__N_166 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_27__7__N_166 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_26__7__N_163 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_26__7__N_163 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_25__7__N_160 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_25__7__N_160 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_24__7__N_157 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_24__7__N_157 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_23__7__N_154 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_23__7__N_154 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_22__7__N_151 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_22__7__N_151 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_21__7__N_148 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_21__7__N_148 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_63__7__N_274 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_63__7__N_274 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_20__7__N_145 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_20__7__N_145 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_19__7__N_142 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_19__7__N_142 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_18__7__N_139 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_18__7__N_139 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_17__7__N_136 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_17__7__N_136 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_16__7__N_133 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_16__7__N_133 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_15__7__N_130 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_15__7__N_130 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_14__7__N_127 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_14__7__N_127 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_13__7__N_124 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_13__7__N_124 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_12__7__N_121 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_12__7__N_121 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_11__7__N_118 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_11__7__N_118 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_10__7__N_115 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_10__7__N_115 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_9__7__N_112 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_9__7__N_112 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_8__7__N_109 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_8__7__N_109 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_7__7__N_106 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_7__7__N_106 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_6__7__N_103 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_6__7__N_103 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_5__7__N_100 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_5__7__N_100 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_4__7__N_97 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_4__7__N_97 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_3__7__N_94 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_3__7__N_94 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_2__7__N_91 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_2__7__N_91 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_1__7__N_88 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_1__7__N_88 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_0__7__N_83 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_0__7__N_83 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[0] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[1] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1453;
    wire [7:0]\mem[62] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[63] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1778, n1391;
    wire [7:0]\mem[2] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[3] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1392;
    wire [7:0]\mem[4] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[5] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1393;
    wire [7:0]\mem[6] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[7] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1394, n1701, n1702, n1717;
    wire [7:0]\mem[32] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[33] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1577, n1703, n1704, n1718, n1608, n1609, n1624;
    wire [7:0]\mem[61] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[34] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[35] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1578;
    wire [7:0]\mem[8] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[9] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1395;
    wire [7:0]\mem[10] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[11] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1396;
    wire [7:0]\mem[12] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[13] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1397, n1610, n1611, n1625;
    wire [7:0]\mem[14] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[15] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1398;
    wire [7:0]\mem[16] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[17] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1399;
    wire [7:0]\mem[18] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[19] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1400;
    wire [7:0]\mem[42] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[43] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1644, n1705, n1706, n1719, n1707, n1708, n1720, n1612, 
        n1613, n1626;
    wire [7:0]\mem[40] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[41] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1643, n1614, n1615, n1627, n1709, n1710, n1721, n1462, 
        n1616, n1617, n1628;
    wire [7:0]\mem[36] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[37] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1579;
    wire [7:0]\mem[38] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[39] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1580, n1581, n1642, n1582;
    wire [7:0]\mem[20] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[21] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1401;
    wire [7:0]\mem[22] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[23] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1402;
    wire [7:0]\mem[24] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[25] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1403;
    wire [7:0]\mem[26] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[27] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1404;
    wire [7:0]\mem[28] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[29] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1405;
    wire [7:0]\mem[30] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[31] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1406, n1641;
    wire [7:0]\mem[44] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[45] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1583;
    wire [7:0]\mem[46] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[47] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1584, n1517, n1516, n1515, n1764, n1763, n1732, n1733, 
        n1748, n1311, n1310, n1654;
    wire [7:0]\mem[60] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1653, n1522;
    wire [7:0]\mem[59] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[58] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[57] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[56] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[55] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[54] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[53] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[52] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[51] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[50] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[49] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[48] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1521, n1769, n1770, n1782, n1640, n1618, n1619, n1629, 
        n1520, n1767, n1519, n1766, n1530, n1765, n1529, n1587, 
        n1588, n1598, n1461, n1473, n1422, n1423, n1438, n1463, 
        n1464, n1474, n1528, n1455, n1456, n1470, n1652, n1525, 
        n1526, n1536, n1620, n1621, n1630, n1622, n1623, n1631, 
        n1465, n1466, n1475, n1651, n1527, n1537, n1499, n1711, 
        n1712, n1722, n1498, n1497, n1496, n1457, n1458, n1471, 
        n1424, n1425, n1439, n1467, n1468, n1476, n1650, n1649, 
        n1495, n1713, n1714, n1723, n1494, n1715, n1716, n1724, 
        n1493, n1492, n1298, n1299, n1314;
    wire [7:0]data_7__N_66;
    
    wire n1648, n1312, n1313, n1321, n1647, n1491, n1490, n1300, 
        n1301, n1315, n1591, n1592, n1600, n1543, n1544, n1545, 
        n1574, n1575, n1576, n1512, n1513, n1514, n1605, n1606, 
        n1607, n1481, n1482, n1483, n1636, n1637, n1638, n1450, 
        n1451, n1452, n1667, n1668, n1669, n1419, n1420, n1421, 
        n1698, n1699, n1700, n1388, n1389, n1390, n1489, n1302, 
        n1303, n1316, n1729, n1730, n1731, n1357, n1358, n1359, 
        n1760, n1761, n1762, n1326, n1327, n1328, n1791, n1792, 
        n1793, n1329, n1330, n1331, n1332, n1488, n1333, n1334, 
        n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
        n1343, n1344, n1736, n1737, n1670, n1671, n1672, n1673, 
        n1304, n1305, n1317, n1546, n1547, n1674, n1675, n1738, 
        n1739, n1771, n1772, n1548, n1734, n1735, n1749, n1549, 
        n1550, n1896, n1551, n1676, n1677, n1552, n1553, n1554, 
        n1555, n1678, n1679, n1740, n1741, n1426, n1427, n1440, 
        n1360, n1361, n1556, n1557, n1362, n1363, n1558, n1559, 
        n1680, n1681, n1364, n1365, n1366, n1367, n1560, n1561, 
        n1682, n1683, n1742, n1743, n1368, n1369, n1370, n1371, 
        n1372, n1373, n1374, n1428, n1429, n1441, n1375, n1684, 
        n1685, n1744, n1745, n1773, n1774, n1306, n1307, n1746, 
        n1747, n1775, n1776, n1777, n1639, n1430, n1431, n1442, 
        n1646, n1432, n1433, n1443, n1437, n1645, n1436, n1487, 
        n1486, n1434, n1435, n1444, n1485, n1445, n1589, n1590, 
        n1599, n1484, n1655, n1459, n1460, n1472, n1656, n1657, 
        n1500, n1501, n1658, n1308, n1309, n1319, n1502, n1518, 
        n1585, n1524, n1523, n1586, n1503, n1659, n1504, n1454, 
        n1768, n1505, n1660, n1506, n1507, n1661, n1780, n1538, 
        n1533, n1781, n1534, n1535, n1662, n1320, n1779, n1531, 
        n1532, n1469, n1597, n1596, n1414, n1413, n1412, n1595, 
        n1594, n1411, n1410, n1409, n1593, n1408, n1407, n1786, 
        n1785, n1755, n1318, n1784, n1754, n1693, n1383, n1382, 
        n1381, n1380, n1753, n1692, n1569, n1379, n1378, n1691, 
        n1568, n1377, n1567, n1376, n1752, n1690, n1566, n1565, 
        n1689, n1564, n1563, n1783, n1751, n1688, n1562, n1687, 
        n1686, n1750, n1352, n1351, n1350, n1349, n1348, n1347, 
        n1346, n1345, n1542, n1541, n1540, n1539, n1666, n1665, 
        n1664, n1663, n1511, n1510, n1509, n1508, n1449, n1448, 
        n1447, n1446, n1325, n1728, n1727, n1324, n1323, n1322, 
        n1726, n1725, n1635, n1634, n1633, n1632, n1790, n1789, 
        n1477, n1478, n1479, n1480, n1604, n1603, n1602, n1601, 
        n1788, n1787, n1418, n1417, n1416, n1415, n1759, n1758, 
        n1757, n1387, n1386, n1385, n1756, n1697, n1696, n1695, 
        n1694, n1573, n1572, n1571, n1384, n1570, n1356, n1355, 
        n1354, n1353;
    
    LUT4 i1383_3_lut (.A(\mem[0] [2]), .B(\mem[1] [2]), .C(address[0]), 
         .Z(n1453)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1383_3_lut.init = 16'hcaca;
    LUT4 i1708_3_lut (.A(\mem[62] [1]), .B(\mem[63] [1]), .C(address[0]), 
         .Z(n1778)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1708_3_lut.init = 16'hcaca;
    LUT4 i1321_3_lut (.A(\mem[0] [3]), .B(\mem[1] [3]), .C(address[0]), 
         .Z(n1391)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1321_3_lut.init = 16'hcaca;
    LUT4 i1322_3_lut (.A(\mem[2] [3]), .B(\mem[3] [3]), .C(address[0]), 
         .Z(n1392)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1322_3_lut.init = 16'hcaca;
    LUT4 i1323_3_lut (.A(\mem[4] [3]), .B(\mem[5] [3]), .C(address[0]), 
         .Z(n1393)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1323_3_lut.init = 16'hcaca;
    LUT4 i1324_3_lut (.A(\mem[6] [3]), .B(\mem[7] [3]), .C(address[0]), 
         .Z(n1394)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1324_3_lut.init = 16'hcaca;
    PFUMX i1647 (.BLUT(n1701), .ALUT(n1702), .C0(address[1]), .Z(n1717));
    LUT4 i1507_3_lut (.A(\mem[32] [0]), .B(\mem[33] [0]), .C(address[0]), 
         .Z(n1577)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1507_3_lut.init = 16'hcaca;
    FD1S1AY data_7__I_0_5187_i1 (.D(data[0]), .CK(mem_62__7__N_271), .Q(\mem[62] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i1.GSR = "DISABLED";
    PFUMX i1648 (.BLUT(n1703), .ALUT(n1704), .C0(address[1]), .Z(n1718));
    PFUMX i1554 (.BLUT(n1608), .ALUT(n1609), .C0(address[1]), .Z(n1624));
    FD1S1A data_7__I_0_5184_i1 (.D(data[0]), .CK(mem_61__7__N_268), .Q(\mem[61] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i1.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut (.A(address[4]), .B(address[5]), .C(address[3]), 
         .Z(n1290)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut.init = 16'hefef;
    LUT4 i1508_3_lut (.A(\mem[34] [0]), .B(\mem[35] [0]), .C(address[0]), 
         .Z(n1578)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1508_3_lut.init = 16'hcaca;
    LUT4 i1325_3_lut (.A(\mem[8] [3]), .B(\mem[9] [3]), .C(address[0]), 
         .Z(n1395)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1325_3_lut.init = 16'hcaca;
    LUT4 i1326_3_lut (.A(\mem[10] [3]), .B(\mem[11] [3]), .C(address[0]), 
         .Z(n1396)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1326_3_lut.init = 16'hcaca;
    LUT4 i1327_3_lut (.A(\mem[12] [3]), .B(\mem[13] [3]), .C(address[0]), 
         .Z(n1397)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1327_3_lut.init = 16'hcaca;
    PFUMX i1555 (.BLUT(n1610), .ALUT(n1611), .C0(address[1]), .Z(n1625));
    LUT4 i1328_3_lut (.A(\mem[14] [3]), .B(\mem[15] [3]), .C(address[0]), 
         .Z(n1398)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1328_3_lut.init = 16'hcaca;
    LUT4 i1329_3_lut (.A(\mem[16] [3]), .B(\mem[17] [3]), .C(address[0]), 
         .Z(n1399)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1329_3_lut.init = 16'hcaca;
    LUT4 i1330_3_lut (.A(\mem[18] [3]), .B(\mem[19] [3]), .C(address[0]), 
         .Z(n1400)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1330_3_lut.init = 16'hcaca;
    LUT4 i1574_3_lut (.A(\mem[42] [6]), .B(\mem[43] [6]), .C(address[0]), 
         .Z(n1644)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1574_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_63 (.A(address[4]), .B(address[5]), .C(address[3]), 
         .Z(n1289)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_adj_63.init = 16'hfefe;
    PFUMX i1649 (.BLUT(n1705), .ALUT(n1706), .C0(address[1]), .Z(n1719));
    PFUMX i1650 (.BLUT(n1707), .ALUT(n1708), .C0(address[1]), .Z(n1720));
    PFUMX i1556 (.BLUT(n1612), .ALUT(n1613), .C0(address[1]), .Z(n1626));
    LUT4 i1573_3_lut (.A(\mem[40] [6]), .B(\mem[41] [6]), .C(address[0]), 
         .Z(n1643)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1573_3_lut.init = 16'hcaca;
    PFUMX i1557 (.BLUT(n1614), .ALUT(n1615), .C0(address[1]), .Z(n1627));
    PFUMX i1651 (.BLUT(n1709), .ALUT(n1710), .C0(address[1]), .Z(n1721));
    LUT4 i1392_3_lut (.A(\mem[18] [2]), .B(\mem[19] [2]), .C(address[0]), 
         .Z(n1462)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1392_3_lut.init = 16'hcaca;
    PFUMX i1558 (.BLUT(n1616), .ALUT(n1617), .C0(address[1]), .Z(n1628));
    LUT4 i1509_3_lut (.A(\mem[36] [0]), .B(\mem[37] [0]), .C(address[0]), 
         .Z(n1579)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1509_3_lut.init = 16'hcaca;
    LUT4 i1510_3_lut (.A(\mem[38] [0]), .B(\mem[39] [0]), .C(address[0]), 
         .Z(n1580)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1510_3_lut.init = 16'hcaca;
    LUT4 i1511_3_lut (.A(\mem[40] [0]), .B(\mem[41] [0]), .C(address[0]), 
         .Z(n1581)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1511_3_lut.init = 16'hcaca;
    LUT4 i1572_3_lut (.A(\mem[38] [6]), .B(\mem[39] [6]), .C(address[0]), 
         .Z(n1642)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1572_3_lut.init = 16'hcaca;
    LUT4 i1512_3_lut (.A(\mem[42] [0]), .B(\mem[43] [0]), .C(address[0]), 
         .Z(n1582)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1512_3_lut.init = 16'hcaca;
    LUT4 i1331_3_lut (.A(\mem[20] [3]), .B(\mem[21] [3]), .C(address[0]), 
         .Z(n1401)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1331_3_lut.init = 16'hcaca;
    LUT4 i1332_3_lut (.A(\mem[22] [3]), .B(\mem[23] [3]), .C(address[0]), 
         .Z(n1402)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1332_3_lut.init = 16'hcaca;
    LUT4 i1333_3_lut (.A(\mem[24] [3]), .B(\mem[25] [3]), .C(address[0]), 
         .Z(n1403)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1333_3_lut.init = 16'hcaca;
    LUT4 i1334_3_lut (.A(\mem[26] [3]), .B(\mem[27] [3]), .C(address[0]), 
         .Z(n1404)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1334_3_lut.init = 16'hcaca;
    LUT4 i1335_3_lut (.A(\mem[28] [3]), .B(\mem[29] [3]), .C(address[0]), 
         .Z(n1405)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1335_3_lut.init = 16'hcaca;
    LUT4 i1336_3_lut (.A(\mem[30] [3]), .B(\mem[31] [3]), .C(address[0]), 
         .Z(n1406)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1336_3_lut.init = 16'hcaca;
    LUT4 i1571_3_lut (.A(\mem[36] [6]), .B(\mem[37] [6]), .C(address[0]), 
         .Z(n1641)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1571_3_lut.init = 16'hcaca;
    LUT4 i1513_3_lut (.A(\mem[44] [0]), .B(\mem[45] [0]), .C(address[0]), 
         .Z(n1583)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1513_3_lut.init = 16'hcaca;
    LUT4 i1514_3_lut (.A(\mem[46] [0]), .B(\mem[47] [0]), .C(address[0]), 
         .Z(n1584)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1514_3_lut.init = 16'hcaca;
    LUT4 i1447_3_lut (.A(\mem[4] [7]), .B(\mem[5] [7]), .C(address[0]), 
         .Z(n1517)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1447_3_lut.init = 16'hcaca;
    LUT4 i1446_3_lut (.A(\mem[2] [7]), .B(\mem[3] [7]), .C(address[0]), 
         .Z(n1516)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1446_3_lut.init = 16'hcaca;
    LUT4 i1445_3_lut (.A(\mem[0] [7]), .B(\mem[1] [7]), .C(address[0]), 
         .Z(n1515)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1445_3_lut.init = 16'hcaca;
    LUT4 i1694_3_lut (.A(\mem[34] [1]), .B(\mem[35] [1]), .C(address[0]), 
         .Z(n1764)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1694_3_lut.init = 16'hcaca;
    LUT4 i1693_3_lut (.A(\mem[32] [1]), .B(\mem[33] [1]), .C(address[0]), 
         .Z(n1763)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1693_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_64 (.A(address[3]), .B(address[5]), .C(address[4]), 
         .Z(n1283)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_adj_64.init = 16'hbfbf;
    PFUMX i1678 (.BLUT(n1732), .ALUT(n1733), .C0(address[1]), .Z(n1748));
    LUT4 i1241_3_lut (.A(\mem[26] [1]), .B(\mem[27] [1]), .C(address[0]), 
         .Z(n1311)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1241_3_lut.init = 16'hcaca;
    LUT4 i1240_3_lut (.A(\mem[24] [1]), .B(\mem[25] [1]), .C(address[0]), 
         .Z(n1310)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1240_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_65 (.A(address[3]), .B(address[5]), .C(address[4]), 
         .Z(n1284)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_adj_65.init = 16'hfbfb;
    LUT4 i1584_3_lut (.A(\mem[62] [6]), .B(\mem[63] [6]), .C(address[0]), 
         .Z(n1654)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1584_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_66 (.A(address[2]), .B(address[0]), .C(address[1]), 
         .Z(n1293)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_adj_66.init = 16'hbfbf;
    LUT4 i1583_3_lut (.A(\mem[60] [6]), .B(\mem[61] [6]), .C(address[0]), 
         .Z(n1653)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1583_3_lut.init = 16'hcaca;
    LUT4 i1452_3_lut (.A(\mem[14] [7]), .B(\mem[15] [7]), .C(address[0]), 
         .Z(n1522)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1452_3_lut.init = 16'hcaca;
    FD1S1A data_7__I_0_5181_i1 (.D(data[0]), .CK(mem_60__7__N_265), .Q(\mem[60] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i1 (.D(data[0]), .CK(mem_59__7__N_262), .Q(\mem[59] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i1 (.D(data[0]), .CK(mem_58__7__N_259), .Q(\mem[58] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i1 (.D(data[0]), .CK(mem_57__7__N_256), .Q(\mem[57] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i1 (.D(data[0]), .CK(mem_56__7__N_253), .Q(\mem[56] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i1 (.D(data[0]), .CK(mem_55__7__N_250), .Q(\mem[55] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i1 (.D(data[0]), .CK(mem_54__7__N_247), .Q(\mem[54] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i1 (.D(data[0]), .CK(mem_53__7__N_244), .Q(\mem[53] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i1 (.D(data[0]), .CK(mem_52__7__N_241), .Q(\mem[52] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i1 (.D(data[0]), .CK(mem_51__7__N_238), .Q(\mem[51] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i1 (.D(data[0]), .CK(mem_50__7__N_235), .Q(\mem[50] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i1 (.D(data[0]), .CK(mem_49__7__N_232), .Q(\mem[49] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i1 (.D(data[0]), .CK(mem_48__7__N_229), .Q(\mem[48] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i1 (.D(data[0]), .CK(mem_47__7__N_226), .Q(\mem[47] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i1 (.D(data[0]), .CK(mem_46__7__N_223), .Q(\mem[46] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i1 (.D(data[0]), .CK(mem_45__7__N_220), .Q(\mem[45] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i1 (.D(data[0]), .CK(mem_44__7__N_217), .Q(\mem[44] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i1 (.D(data[0]), .CK(mem_43__7__N_214), .Q(\mem[43] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i1 (.D(data[0]), .CK(mem_42__7__N_211), .Q(\mem[42] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i1 (.D(data[0]), .CK(mem_41__7__N_208), .Q(\mem[41] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i1 (.D(data[0]), .CK(mem_40__7__N_205), .Q(\mem[40] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i1 (.D(data[0]), .CK(mem_39__7__N_202), .Q(\mem[39] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i1 (.D(data[0]), .CK(mem_38__7__N_199), .Q(\mem[38] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i1 (.D(data[0]), .CK(mem_37__7__N_196), .Q(\mem[37] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i1 (.D(data[0]), .CK(mem_36__7__N_193), .Q(\mem[36] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i1 (.D(data[0]), .CK(mem_35__7__N_190), .Q(\mem[35] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i1 (.D(data[0]), .CK(mem_34__7__N_187), .Q(\mem[34] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i1 (.D(data[0]), .CK(mem_33__7__N_184), .Q(\mem[33] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i1 (.D(data[0]), .CK(mem_32__7__N_181), .Q(\mem[32] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i1 (.D(data[0]), .CK(mem_31__7__N_178), .Q(\mem[31] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i1 (.D(data[0]), .CK(mem_30__7__N_175), .Q(\mem[30] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i1 (.D(data[0]), .CK(mem_29__7__N_172), .Q(\mem[29] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i1 (.D(data[0]), .CK(mem_28__7__N_169), .Q(\mem[28] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i1 (.D(data[0]), .CK(mem_27__7__N_166), .Q(\mem[27] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i1 (.D(data[0]), .CK(mem_26__7__N_163), .Q(\mem[26] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i1 (.D(data[0]), .CK(mem_25__7__N_160), .Q(\mem[25] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i1.GSR = "DISABLED";
    LUT4 i1451_3_lut (.A(\mem[12] [7]), .B(\mem[13] [7]), .C(address[0]), 
         .Z(n1521)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1451_3_lut.init = 16'hcaca;
    PFUMX i1712 (.BLUT(n1769), .ALUT(n1770), .C0(address[1]), .Z(n1782));
    FD1S1A data_7__I_0_5073_i1 (.D(data[0]), .CK(mem_24__7__N_157), .Q(\mem[24] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i1 (.D(data[0]), .CK(mem_23__7__N_154), .Q(\mem[23] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i1 (.D(data[0]), .CK(mem_22__7__N_151), .Q(\mem[22] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i1 (.D(data[0]), .CK(mem_21__7__N_148), .Q(\mem[21] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i1.GSR = "DISABLED";
    FD1S1AY data_7__I_0_i1 (.D(data[0]), .CK(mem_63__7__N_274), .Q(\mem[63] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i1.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5061_i1 (.D(data[0]), .CK(mem_20__7__N_145), .Q(\mem[20] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i1.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5058_i1 (.D(data[0]), .CK(mem_19__7__N_142), .Q(\mem[19] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i1.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5055_i1 (.D(data[0]), .CK(mem_18__7__N_139), .Q(\mem[18] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i1.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5052_i1 (.D(data[0]), .CK(mem_17__7__N_136), .Q(\mem[17] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i1 (.D(data[0]), .CK(mem_16__7__N_133), .Q(\mem[16] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i1.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5046_i1 (.D(data[0]), .CK(mem_15__7__N_130), .Q(\mem[15] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i1.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5043_i1 (.D(data[0]), .CK(mem_14__7__N_127), .Q(\mem[14] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5040_i1 (.D(data[0]), .CK(mem_13__7__N_124), .Q(\mem[13] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i1.GSR = "DISABLED";
    LUT4 i1570_3_lut (.A(\mem[34] [6]), .B(\mem[35] [6]), .C(address[0]), 
         .Z(n1640)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1570_3_lut.init = 16'hcaca;
    FD1S1AY data_7__I_0_5037_i1 (.D(data[0]), .CK(mem_12__7__N_121), .Q(\mem[12] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i1 (.D(data[0]), .CK(mem_11__7__N_118), .Q(\mem[11] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5031_i1 (.D(data[0]), .CK(mem_10__7__N_115), .Q(\mem[10] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5028_i1 (.D(data[0]), .CK(mem_9__7__N_112), .Q(\mem[9] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i1.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5025_i1 (.D(data[0]), .CK(mem_8__7__N_109), .Q(\mem[8] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5022_i1 (.D(data[0]), .CK(mem_7__7__N_106), .Q(\mem[7] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i1.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5019_i1 (.D(data[0]), .CK(mem_6__7__N_103), .Q(\mem[6] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i1.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5016_i1 (.D(data[0]), .CK(mem_5__7__N_100), .Q(\mem[5] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5013_i1 (.D(data[0]), .CK(mem_4__7__N_97), .Q(\mem[4] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i1.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5010_i1 (.D(data[0]), .CK(mem_3__7__N_94), .Q(\mem[3] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i1.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5007_i1 (.D(data[0]), .CK(mem_2__7__N_91), .Q(\mem[2] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5004_i1 (.D(data[0]), .CK(mem_1__7__N_88), .Q(\mem[1] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5002_i1 (.D(data[0]), .CK(mem_0__7__N_83), .Q(\mem[0] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i1.GSR = "DISABLED";
    PFUMX i1559 (.BLUT(n1618), .ALUT(n1619), .C0(address[1]), .Z(n1629));
    LUT4 i1450_3_lut (.A(\mem[10] [7]), .B(\mem[11] [7]), .C(address[0]), 
         .Z(n1520)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1450_3_lut.init = 16'hcaca;
    FD1S1AY data_7__I_0_5002_i2 (.D(data[1]), .CK(mem_0__7__N_83), .Q(\mem[0] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5002_i3 (.D(data[2]), .CK(mem_0__7__N_83), .Q(\mem[0] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i3.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5002_i4 (.D(data[3]), .CK(mem_0__7__N_83), .Q(\mem[0] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i4.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5002_i5 (.D(data[4]), .CK(mem_0__7__N_83), .Q(\mem[0] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i5.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5002_i6 (.D(data[5]), .CK(mem_0__7__N_83), .Q(\mem[0] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5002_i7 (.D(data[6]), .CK(mem_0__7__N_83), .Q(\mem[0] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5002_i8 (.D(data[7]), .CK(mem_0__7__N_83), .Q(\mem[0] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5004_i2 (.D(data[1]), .CK(mem_1__7__N_88), .Q(\mem[1] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5004_i3 (.D(data[2]), .CK(mem_1__7__N_88), .Q(\mem[1] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5004_i4 (.D(data[3]), .CK(mem_1__7__N_88), .Q(\mem[1] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i4.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5004_i5 (.D(data[4]), .CK(mem_1__7__N_88), .Q(\mem[1] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5004_i6 (.D(data[5]), .CK(mem_1__7__N_88), .Q(\mem[1] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5004_i7 (.D(data[6]), .CK(mem_1__7__N_88), .Q(\mem[1] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5004_i8 (.D(data[7]), .CK(mem_1__7__N_88), .Q(\mem[1] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i8.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5007_i2 (.D(data[1]), .CK(mem_2__7__N_91), .Q(\mem[2] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5007_i3 (.D(data[2]), .CK(mem_2__7__N_91), .Q(\mem[2] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i3.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5007_i4 (.D(data[3]), .CK(mem_2__7__N_91), .Q(\mem[2] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i4.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5007_i5 (.D(data[4]), .CK(mem_2__7__N_91), .Q(\mem[2] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i5.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5007_i6 (.D(data[5]), .CK(mem_2__7__N_91), .Q(\mem[2] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i6.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5007_i7 (.D(data[6]), .CK(mem_2__7__N_91), .Q(\mem[2] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5007_i8 (.D(data[7]), .CK(mem_2__7__N_91), .Q(\mem[2] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5010_i2 (.D(data[1]), .CK(mem_3__7__N_94), .Q(\mem[3] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5010_i3 (.D(data[2]), .CK(mem_3__7__N_94), .Q(\mem[3] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5010_i4 (.D(data[3]), .CK(mem_3__7__N_94), .Q(\mem[3] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i4.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5010_i5 (.D(data[4]), .CK(mem_3__7__N_94), .Q(\mem[3] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5010_i6 (.D(data[5]), .CK(mem_3__7__N_94), .Q(\mem[3] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5010_i7 (.D(data[6]), .CK(mem_3__7__N_94), .Q(\mem[3] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i7.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5010_i8 (.D(data[7]), .CK(mem_3__7__N_94), .Q(\mem[3] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i8.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5013_i2 (.D(data[1]), .CK(mem_4__7__N_97), .Q(\mem[4] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5013_i3 (.D(data[2]), .CK(mem_4__7__N_97), .Q(\mem[4] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i3.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5013_i4 (.D(data[3]), .CK(mem_4__7__N_97), .Q(\mem[4] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i4.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5013_i5 (.D(data[4]), .CK(mem_4__7__N_97), .Q(\mem[4] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i5.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5013_i6 (.D(data[5]), .CK(mem_4__7__N_97), .Q(\mem[4] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5013_i7 (.D(data[6]), .CK(mem_4__7__N_97), .Q(\mem[4] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5013_i8 (.D(data[7]), .CK(mem_4__7__N_97), .Q(\mem[4] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5016_i2 (.D(data[1]), .CK(mem_5__7__N_100), .Q(\mem[5] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5016_i3 (.D(data[2]), .CK(mem_5__7__N_100), .Q(\mem[5] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5016_i4 (.D(data[3]), .CK(mem_5__7__N_100), .Q(\mem[5] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i4.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5016_i5 (.D(data[4]), .CK(mem_5__7__N_100), .Q(\mem[5] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5016_i6 (.D(data[5]), .CK(mem_5__7__N_100), .Q(\mem[5] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i6.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5016_i7 (.D(data[6]), .CK(mem_5__7__N_100), .Q(\mem[5] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5016_i8 (.D(data[7]), .CK(mem_5__7__N_100), .Q(\mem[5] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i8.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5019_i2 (.D(data[1]), .CK(mem_6__7__N_103), .Q(\mem[6] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5019_i3 (.D(data[2]), .CK(mem_6__7__N_103), .Q(\mem[6] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5019_i4 (.D(data[3]), .CK(mem_6__7__N_103), .Q(\mem[6] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i4.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5019_i5 (.D(data[4]), .CK(mem_6__7__N_103), .Q(\mem[6] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5019_i6 (.D(data[5]), .CK(mem_6__7__N_103), .Q(\mem[6] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i6.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5019_i7 (.D(data[6]), .CK(mem_6__7__N_103), .Q(\mem[6] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5019_i8 (.D(data[7]), .CK(mem_6__7__N_103), .Q(\mem[6] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5022_i2 (.D(data[1]), .CK(mem_7__7__N_106), .Q(\mem[7] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5022_i3 (.D(data[2]), .CK(mem_7__7__N_106), .Q(\mem[7] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i3.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5022_i4 (.D(data[3]), .CK(mem_7__7__N_106), .Q(\mem[7] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5022_i5 (.D(data[4]), .CK(mem_7__7__N_106), .Q(\mem[7] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5022_i6 (.D(data[5]), .CK(mem_7__7__N_106), .Q(\mem[7] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i6.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5022_i7 (.D(data[6]), .CK(mem_7__7__N_106), .Q(\mem[7] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i7.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5022_i8 (.D(data[7]), .CK(mem_7__7__N_106), .Q(\mem[7] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i8.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5025_i2 (.D(data[1]), .CK(mem_8__7__N_109), .Q(\mem[8] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5025_i3 (.D(data[2]), .CK(mem_8__7__N_109), .Q(\mem[8] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5025_i4 (.D(data[3]), .CK(mem_8__7__N_109), .Q(\mem[8] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i4.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5025_i5 (.D(data[4]), .CK(mem_8__7__N_109), .Q(\mem[8] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5025_i6 (.D(data[5]), .CK(mem_8__7__N_109), .Q(\mem[8] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5025_i7 (.D(data[6]), .CK(mem_8__7__N_109), .Q(\mem[8] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i7.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5025_i8 (.D(data[7]), .CK(mem_8__7__N_109), .Q(\mem[8] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i8.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5028_i2 (.D(data[1]), .CK(mem_9__7__N_112), .Q(\mem[9] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5028_i3 (.D(data[2]), .CK(mem_9__7__N_112), .Q(\mem[9] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i3.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5028_i4 (.D(data[3]), .CK(mem_9__7__N_112), .Q(\mem[9] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i4.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5028_i5 (.D(data[4]), .CK(mem_9__7__N_112), .Q(\mem[9] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i5.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5028_i6 (.D(data[5]), .CK(mem_9__7__N_112), .Q(\mem[9] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i6.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5028_i7 (.D(data[6]), .CK(mem_9__7__N_112), .Q(\mem[9] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5028_i8 (.D(data[7]), .CK(mem_9__7__N_112), .Q(\mem[9] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i8.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5031_i2 (.D(data[1]), .CK(mem_10__7__N_115), .Q(\mem[10] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5031_i3 (.D(data[2]), .CK(mem_10__7__N_115), .Q(\mem[10] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i3.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5031_i4 (.D(data[3]), .CK(mem_10__7__N_115), .Q(\mem[10] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5031_i5 (.D(data[4]), .CK(mem_10__7__N_115), .Q(\mem[10] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5031_i6 (.D(data[5]), .CK(mem_10__7__N_115), .Q(\mem[10] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i6.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5031_i7 (.D(data[6]), .CK(mem_10__7__N_115), .Q(\mem[10] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i7.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5031_i8 (.D(data[7]), .CK(mem_10__7__N_115), .Q(\mem[10] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i2 (.D(data[1]), .CK(mem_11__7__N_118), .Q(\mem[11] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5034_i3 (.D(data[2]), .CK(mem_11__7__N_118), .Q(\mem[11] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i4 (.D(data[3]), .CK(mem_11__7__N_118), .Q(\mem[11] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i5 (.D(data[4]), .CK(mem_11__7__N_118), .Q(\mem[11] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i6 (.D(data[5]), .CK(mem_11__7__N_118), .Q(\mem[11] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i6.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5034_i7 (.D(data[6]), .CK(mem_11__7__N_118), .Q(\mem[11] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i7.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5034_i8 (.D(data[7]), .CK(mem_11__7__N_118), .Q(\mem[11] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5037_i2 (.D(data[1]), .CK(mem_12__7__N_121), .Q(\mem[12] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5037_i3 (.D(data[2]), .CK(mem_12__7__N_121), .Q(\mem[12] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5037_i4 (.D(data[3]), .CK(mem_12__7__N_121), .Q(\mem[12] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i4.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5037_i5 (.D(data[4]), .CK(mem_12__7__N_121), .Q(\mem[12] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5037_i6 (.D(data[5]), .CK(mem_12__7__N_121), .Q(\mem[12] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5037_i7 (.D(data[6]), .CK(mem_12__7__N_121), .Q(\mem[12] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i7.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5037_i8 (.D(data[7]), .CK(mem_12__7__N_121), .Q(\mem[12] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i8.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5040_i2 (.D(data[1]), .CK(mem_13__7__N_124), .Q(\mem[13] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5040_i3 (.D(data[2]), .CK(mem_13__7__N_124), .Q(\mem[13] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5040_i4 (.D(data[3]), .CK(mem_13__7__N_124), .Q(\mem[13] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5040_i5 (.D(data[4]), .CK(mem_13__7__N_124), .Q(\mem[13] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5040_i6 (.D(data[5]), .CK(mem_13__7__N_124), .Q(\mem[13] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i6.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5040_i7 (.D(data[6]), .CK(mem_13__7__N_124), .Q(\mem[13] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i7.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5040_i8 (.D(data[7]), .CK(mem_13__7__N_124), .Q(\mem[13] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5043_i2 (.D(data[1]), .CK(mem_14__7__N_127), .Q(\mem[14] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5043_i3 (.D(data[2]), .CK(mem_14__7__N_127), .Q(\mem[14] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5043_i4 (.D(data[3]), .CK(mem_14__7__N_127), .Q(\mem[14] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i4.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5043_i5 (.D(data[4]), .CK(mem_14__7__N_127), .Q(\mem[14] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5043_i6 (.D(data[5]), .CK(mem_14__7__N_127), .Q(\mem[14] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i6.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5043_i7 (.D(data[6]), .CK(mem_14__7__N_127), .Q(\mem[14] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5043_i8 (.D(data[7]), .CK(mem_14__7__N_127), .Q(\mem[14] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5046_i2 (.D(data[1]), .CK(mem_15__7__N_130), .Q(\mem[15] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5046_i3 (.D(data[2]), .CK(mem_15__7__N_130), .Q(\mem[15] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i3.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5046_i4 (.D(data[3]), .CK(mem_15__7__N_130), .Q(\mem[15] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i4.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5046_i5 (.D(data[4]), .CK(mem_15__7__N_130), .Q(\mem[15] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i5.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5046_i6 (.D(data[5]), .CK(mem_15__7__N_130), .Q(\mem[15] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5046_i7 (.D(data[6]), .CK(mem_15__7__N_130), .Q(\mem[15] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5046_i8 (.D(data[7]), .CK(mem_15__7__N_130), .Q(\mem[15] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i2 (.D(data[1]), .CK(mem_16__7__N_133), .Q(\mem[16] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5049_i3 (.D(data[2]), .CK(mem_16__7__N_133), .Q(\mem[16] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i4 (.D(data[3]), .CK(mem_16__7__N_133), .Q(\mem[16] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i4.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5049_i5 (.D(data[4]), .CK(mem_16__7__N_133), .Q(\mem[16] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i6 (.D(data[5]), .CK(mem_16__7__N_133), .Q(\mem[16] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i7 (.D(data[6]), .CK(mem_16__7__N_133), .Q(\mem[16] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i7.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5049_i8 (.D(data[7]), .CK(mem_16__7__N_133), .Q(\mem[16] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5052_i2 (.D(data[1]), .CK(mem_17__7__N_136), .Q(\mem[17] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5052_i3 (.D(data[2]), .CK(mem_17__7__N_136), .Q(\mem[17] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5052_i4 (.D(data[3]), .CK(mem_17__7__N_136), .Q(\mem[17] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i4.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5052_i5 (.D(data[4]), .CK(mem_17__7__N_136), .Q(\mem[17] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5052_i6 (.D(data[5]), .CK(mem_17__7__N_136), .Q(\mem[17] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i6.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5052_i7 (.D(data[6]), .CK(mem_17__7__N_136), .Q(\mem[17] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i7.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5052_i8 (.D(data[7]), .CK(mem_17__7__N_136), .Q(\mem[17] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5055_i2 (.D(data[1]), .CK(mem_18__7__N_139), .Q(\mem[18] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5055_i3 (.D(data[2]), .CK(mem_18__7__N_139), .Q(\mem[18] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5055_i4 (.D(data[3]), .CK(mem_18__7__N_139), .Q(\mem[18] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i4.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5055_i5 (.D(data[4]), .CK(mem_18__7__N_139), .Q(\mem[18] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5055_i6 (.D(data[5]), .CK(mem_18__7__N_139), .Q(\mem[18] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i6.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5055_i7 (.D(data[6]), .CK(mem_18__7__N_139), .Q(\mem[18] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i7.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5055_i8 (.D(data[7]), .CK(mem_18__7__N_139), .Q(\mem[18] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i2 (.D(data[1]), .CK(mem_19__7__N_142), .Q(\mem[19] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5058_i3 (.D(data[2]), .CK(mem_19__7__N_142), .Q(\mem[19] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i4 (.D(data[3]), .CK(mem_19__7__N_142), .Q(\mem[19] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i5 (.D(data[4]), .CK(mem_19__7__N_142), .Q(\mem[19] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i6 (.D(data[5]), .CK(mem_19__7__N_142), .Q(\mem[19] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i7 (.D(data[6]), .CK(mem_19__7__N_142), .Q(\mem[19] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i8 (.D(data[7]), .CK(mem_19__7__N_142), .Q(\mem[19] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i8.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5061_i2 (.D(data[1]), .CK(mem_20__7__N_145), .Q(\mem[20] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5061_i3 (.D(data[2]), .CK(mem_20__7__N_145), .Q(\mem[20] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i3.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5061_i4 (.D(data[3]), .CK(mem_20__7__N_145), .Q(\mem[20] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5061_i5 (.D(data[4]), .CK(mem_20__7__N_145), .Q(\mem[20] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5061_i6 (.D(data[5]), .CK(mem_20__7__N_145), .Q(\mem[20] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5061_i7 (.D(data[6]), .CK(mem_20__7__N_145), .Q(\mem[20] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5061_i8 (.D(data[7]), .CK(mem_20__7__N_145), .Q(\mem[20] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_i2 (.D(data[1]), .CK(mem_63__7__N_274), .Q(\mem[63] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_i3 (.D(data[2]), .CK(mem_63__7__N_274), .Q(\mem[63] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_i4 (.D(data[3]), .CK(mem_63__7__N_274), .Q(\mem[63] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_i5 (.D(data[4]), .CK(mem_63__7__N_274), .Q(\mem[63] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_i6 (.D(data[5]), .CK(mem_63__7__N_274), .Q(\mem[63] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_i7 (.D(data[6]), .CK(mem_63__7__N_274), .Q(\mem[63] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_i8 (.D(data[7]), .CK(mem_63__7__N_274), .Q(\mem[63] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i8.GSR = "DISABLED";
    LUT4 i1697_3_lut (.A(\mem[40] [1]), .B(\mem[41] [1]), .C(address[0]), 
         .Z(n1767)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1697_3_lut.init = 16'hcaca;
    LUT4 i1449_3_lut (.A(\mem[8] [7]), .B(\mem[9] [7]), .C(address[0]), 
         .Z(n1519)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1449_3_lut.init = 16'hcaca;
    LUT4 i1696_3_lut (.A(\mem[38] [1]), .B(\mem[39] [1]), .C(address[0]), 
         .Z(n1766)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1696_3_lut.init = 16'hcaca;
    LUT4 i1460_3_lut (.A(\mem[30] [7]), .B(\mem[31] [7]), .C(address[0]), 
         .Z(n1530)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1460_3_lut.init = 16'hcaca;
    LUT4 i1695_3_lut (.A(\mem[36] [1]), .B(\mem[37] [1]), .C(address[0]), 
         .Z(n1765)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1695_3_lut.init = 16'hcaca;
    FD1S1AY data_7__I_0_5187_i2 (.D(data[1]), .CK(mem_62__7__N_271), .Q(\mem[62] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i2.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_adj_67 (.A(address[2]), .B(address[0]), .C(address[1]), 
         .Z(n1292)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_adj_67.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_adj_68 (.A(address[0]), .B(address[1]), .C(address[2]), 
         .Z(n1296)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_adj_68.init = 16'hefef;
    FD1S1AY data_7__I_0_5187_i3 (.D(data[2]), .CK(mem_62__7__N_271), .Q(\mem[62] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i3.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5187_i4 (.D(data[3]), .CK(mem_62__7__N_271), .Q(\mem[62] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i4.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5187_i5 (.D(data[4]), .CK(mem_62__7__N_271), .Q(\mem[62] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i5.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5187_i6 (.D(data[5]), .CK(mem_62__7__N_271), .Q(\mem[62] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i6.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5187_i7 (.D(data[6]), .CK(mem_62__7__N_271), .Q(\mem[62] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i7.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5187_i8 (.D(data[7]), .CK(mem_62__7__N_271), .Q(\mem[62] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i2 (.D(data[1]), .CK(mem_61__7__N_268), .Q(\mem[61] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i3 (.D(data[2]), .CK(mem_61__7__N_268), .Q(\mem[61] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i4 (.D(data[3]), .CK(mem_61__7__N_268), .Q(\mem[61] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i5 (.D(data[4]), .CK(mem_61__7__N_268), .Q(\mem[61] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i6 (.D(data[5]), .CK(mem_61__7__N_268), .Q(\mem[61] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i7 (.D(data[6]), .CK(mem_61__7__N_268), .Q(\mem[61] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i8 (.D(data[7]), .CK(mem_61__7__N_268), .Q(\mem[61] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i2 (.D(data[1]), .CK(mem_60__7__N_265), .Q(\mem[60] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i3 (.D(data[2]), .CK(mem_60__7__N_265), .Q(\mem[60] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i4 (.D(data[3]), .CK(mem_60__7__N_265), .Q(\mem[60] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i5 (.D(data[4]), .CK(mem_60__7__N_265), .Q(\mem[60] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i6 (.D(data[5]), .CK(mem_60__7__N_265), .Q(\mem[60] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i7 (.D(data[6]), .CK(mem_60__7__N_265), .Q(\mem[60] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i8 (.D(data[7]), .CK(mem_60__7__N_265), .Q(\mem[60] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i2 (.D(data[1]), .CK(mem_59__7__N_262), .Q(\mem[59] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i3 (.D(data[2]), .CK(mem_59__7__N_262), .Q(\mem[59] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i4 (.D(data[3]), .CK(mem_59__7__N_262), .Q(\mem[59] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i5 (.D(data[4]), .CK(mem_59__7__N_262), .Q(\mem[59] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i6 (.D(data[5]), .CK(mem_59__7__N_262), .Q(\mem[59] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i7 (.D(data[6]), .CK(mem_59__7__N_262), .Q(\mem[59] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i8 (.D(data[7]), .CK(mem_59__7__N_262), .Q(\mem[59] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i2 (.D(data[1]), .CK(mem_58__7__N_259), .Q(\mem[58] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i3 (.D(data[2]), .CK(mem_58__7__N_259), .Q(\mem[58] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i4 (.D(data[3]), .CK(mem_58__7__N_259), .Q(\mem[58] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i5 (.D(data[4]), .CK(mem_58__7__N_259), .Q(\mem[58] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i6 (.D(data[5]), .CK(mem_58__7__N_259), .Q(\mem[58] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i7 (.D(data[6]), .CK(mem_58__7__N_259), .Q(\mem[58] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i8 (.D(data[7]), .CK(mem_58__7__N_259), .Q(\mem[58] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i2 (.D(data[1]), .CK(mem_57__7__N_256), .Q(\mem[57] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i3 (.D(data[2]), .CK(mem_57__7__N_256), .Q(\mem[57] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i4 (.D(data[3]), .CK(mem_57__7__N_256), .Q(\mem[57] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i5 (.D(data[4]), .CK(mem_57__7__N_256), .Q(\mem[57] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i6 (.D(data[5]), .CK(mem_57__7__N_256), .Q(\mem[57] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i7 (.D(data[6]), .CK(mem_57__7__N_256), .Q(\mem[57] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i8 (.D(data[7]), .CK(mem_57__7__N_256), .Q(\mem[57] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i2 (.D(data[1]), .CK(mem_56__7__N_253), .Q(\mem[56] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i3 (.D(data[2]), .CK(mem_56__7__N_253), .Q(\mem[56] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i4 (.D(data[3]), .CK(mem_56__7__N_253), .Q(\mem[56] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i5 (.D(data[4]), .CK(mem_56__7__N_253), .Q(\mem[56] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i6 (.D(data[5]), .CK(mem_56__7__N_253), .Q(\mem[56] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i7 (.D(data[6]), .CK(mem_56__7__N_253), .Q(\mem[56] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i8 (.D(data[7]), .CK(mem_56__7__N_253), .Q(\mem[56] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i2 (.D(data[1]), .CK(mem_55__7__N_250), .Q(\mem[55] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i3 (.D(data[2]), .CK(mem_55__7__N_250), .Q(\mem[55] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i4 (.D(data[3]), .CK(mem_55__7__N_250), .Q(\mem[55] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i5 (.D(data[4]), .CK(mem_55__7__N_250), .Q(\mem[55] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i6 (.D(data[5]), .CK(mem_55__7__N_250), .Q(\mem[55] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i7 (.D(data[6]), .CK(mem_55__7__N_250), .Q(\mem[55] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i8 (.D(data[7]), .CK(mem_55__7__N_250), .Q(\mem[55] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i2 (.D(data[1]), .CK(mem_54__7__N_247), .Q(\mem[54] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i3 (.D(data[2]), .CK(mem_54__7__N_247), .Q(\mem[54] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i4 (.D(data[3]), .CK(mem_54__7__N_247), .Q(\mem[54] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i5 (.D(data[4]), .CK(mem_54__7__N_247), .Q(\mem[54] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i6 (.D(data[5]), .CK(mem_54__7__N_247), .Q(\mem[54] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i7 (.D(data[6]), .CK(mem_54__7__N_247), .Q(\mem[54] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i8 (.D(data[7]), .CK(mem_54__7__N_247), .Q(\mem[54] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i2 (.D(data[1]), .CK(mem_53__7__N_244), .Q(\mem[53] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i3 (.D(data[2]), .CK(mem_53__7__N_244), .Q(\mem[53] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i4 (.D(data[3]), .CK(mem_53__7__N_244), .Q(\mem[53] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i5 (.D(data[4]), .CK(mem_53__7__N_244), .Q(\mem[53] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i6 (.D(data[5]), .CK(mem_53__7__N_244), .Q(\mem[53] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i7 (.D(data[6]), .CK(mem_53__7__N_244), .Q(\mem[53] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i8 (.D(data[7]), .CK(mem_53__7__N_244), .Q(\mem[53] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i2 (.D(data[1]), .CK(mem_52__7__N_241), .Q(\mem[52] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i3 (.D(data[2]), .CK(mem_52__7__N_241), .Q(\mem[52] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i4 (.D(data[3]), .CK(mem_52__7__N_241), .Q(\mem[52] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i5 (.D(data[4]), .CK(mem_52__7__N_241), .Q(\mem[52] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i6 (.D(data[5]), .CK(mem_52__7__N_241), .Q(\mem[52] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i7 (.D(data[6]), .CK(mem_52__7__N_241), .Q(\mem[52] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i8 (.D(data[7]), .CK(mem_52__7__N_241), .Q(\mem[52] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i2 (.D(data[1]), .CK(mem_51__7__N_238), .Q(\mem[51] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i3 (.D(data[2]), .CK(mem_51__7__N_238), .Q(\mem[51] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i4 (.D(data[3]), .CK(mem_51__7__N_238), .Q(\mem[51] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i5 (.D(data[4]), .CK(mem_51__7__N_238), .Q(\mem[51] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i6 (.D(data[5]), .CK(mem_51__7__N_238), .Q(\mem[51] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i7 (.D(data[6]), .CK(mem_51__7__N_238), .Q(\mem[51] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i8 (.D(data[7]), .CK(mem_51__7__N_238), .Q(\mem[51] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i2 (.D(data[1]), .CK(mem_50__7__N_235), .Q(\mem[50] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i3 (.D(data[2]), .CK(mem_50__7__N_235), .Q(\mem[50] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i4 (.D(data[3]), .CK(mem_50__7__N_235), .Q(\mem[50] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i5 (.D(data[4]), .CK(mem_50__7__N_235), .Q(\mem[50] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i6 (.D(data[5]), .CK(mem_50__7__N_235), .Q(\mem[50] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i7 (.D(data[6]), .CK(mem_50__7__N_235), .Q(\mem[50] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i8 (.D(data[7]), .CK(mem_50__7__N_235), .Q(\mem[50] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i2 (.D(data[1]), .CK(mem_49__7__N_232), .Q(\mem[49] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i3 (.D(data[2]), .CK(mem_49__7__N_232), .Q(\mem[49] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i4 (.D(data[3]), .CK(mem_49__7__N_232), .Q(\mem[49] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i5 (.D(data[4]), .CK(mem_49__7__N_232), .Q(\mem[49] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i6 (.D(data[5]), .CK(mem_49__7__N_232), .Q(\mem[49] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i7 (.D(data[6]), .CK(mem_49__7__N_232), .Q(\mem[49] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i8 (.D(data[7]), .CK(mem_49__7__N_232), .Q(\mem[49] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i2 (.D(data[1]), .CK(mem_48__7__N_229), .Q(\mem[48] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i3 (.D(data[2]), .CK(mem_48__7__N_229), .Q(\mem[48] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i4 (.D(data[3]), .CK(mem_48__7__N_229), .Q(\mem[48] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i5 (.D(data[4]), .CK(mem_48__7__N_229), .Q(\mem[48] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i6 (.D(data[5]), .CK(mem_48__7__N_229), .Q(\mem[48] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i7 (.D(data[6]), .CK(mem_48__7__N_229), .Q(\mem[48] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i8 (.D(data[7]), .CK(mem_48__7__N_229), .Q(\mem[48] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i2 (.D(data[1]), .CK(mem_47__7__N_226), .Q(\mem[47] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i3 (.D(data[2]), .CK(mem_47__7__N_226), .Q(\mem[47] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i4 (.D(data[3]), .CK(mem_47__7__N_226), .Q(\mem[47] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i5 (.D(data[4]), .CK(mem_47__7__N_226), .Q(\mem[47] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i6 (.D(data[5]), .CK(mem_47__7__N_226), .Q(\mem[47] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i7 (.D(data[6]), .CK(mem_47__7__N_226), .Q(\mem[47] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i8 (.D(data[7]), .CK(mem_47__7__N_226), .Q(\mem[47] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i2 (.D(data[1]), .CK(mem_46__7__N_223), .Q(\mem[46] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i3 (.D(data[2]), .CK(mem_46__7__N_223), .Q(\mem[46] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i4 (.D(data[3]), .CK(mem_46__7__N_223), .Q(\mem[46] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i5 (.D(data[4]), .CK(mem_46__7__N_223), .Q(\mem[46] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i6 (.D(data[5]), .CK(mem_46__7__N_223), .Q(\mem[46] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i7 (.D(data[6]), .CK(mem_46__7__N_223), .Q(\mem[46] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i8 (.D(data[7]), .CK(mem_46__7__N_223), .Q(\mem[46] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i2 (.D(data[1]), .CK(mem_45__7__N_220), .Q(\mem[45] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i3 (.D(data[2]), .CK(mem_45__7__N_220), .Q(\mem[45] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i4 (.D(data[3]), .CK(mem_45__7__N_220), .Q(\mem[45] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i5 (.D(data[4]), .CK(mem_45__7__N_220), .Q(\mem[45] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i6 (.D(data[5]), .CK(mem_45__7__N_220), .Q(\mem[45] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i7 (.D(data[6]), .CK(mem_45__7__N_220), .Q(\mem[45] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i8 (.D(data[7]), .CK(mem_45__7__N_220), .Q(\mem[45] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i2 (.D(data[1]), .CK(mem_44__7__N_217), .Q(\mem[44] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i3 (.D(data[2]), .CK(mem_44__7__N_217), .Q(\mem[44] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i4 (.D(data[3]), .CK(mem_44__7__N_217), .Q(\mem[44] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i5 (.D(data[4]), .CK(mem_44__7__N_217), .Q(\mem[44] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i6 (.D(data[5]), .CK(mem_44__7__N_217), .Q(\mem[44] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i7 (.D(data[6]), .CK(mem_44__7__N_217), .Q(\mem[44] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i8 (.D(data[7]), .CK(mem_44__7__N_217), .Q(\mem[44] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i2 (.D(data[1]), .CK(mem_43__7__N_214), .Q(\mem[43] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i3 (.D(data[2]), .CK(mem_43__7__N_214), .Q(\mem[43] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i4 (.D(data[3]), .CK(mem_43__7__N_214), .Q(\mem[43] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i5 (.D(data[4]), .CK(mem_43__7__N_214), .Q(\mem[43] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i6 (.D(data[5]), .CK(mem_43__7__N_214), .Q(\mem[43] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i7 (.D(data[6]), .CK(mem_43__7__N_214), .Q(\mem[43] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i8 (.D(data[7]), .CK(mem_43__7__N_214), .Q(\mem[43] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i2 (.D(data[1]), .CK(mem_42__7__N_211), .Q(\mem[42] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i3 (.D(data[2]), .CK(mem_42__7__N_211), .Q(\mem[42] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i4 (.D(data[3]), .CK(mem_42__7__N_211), .Q(\mem[42] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i5 (.D(data[4]), .CK(mem_42__7__N_211), .Q(\mem[42] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i6 (.D(data[5]), .CK(mem_42__7__N_211), .Q(\mem[42] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i7 (.D(data[6]), .CK(mem_42__7__N_211), .Q(\mem[42] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i8 (.D(data[7]), .CK(mem_42__7__N_211), .Q(\mem[42] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i2 (.D(data[1]), .CK(mem_41__7__N_208), .Q(\mem[41] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i3 (.D(data[2]), .CK(mem_41__7__N_208), .Q(\mem[41] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i4 (.D(data[3]), .CK(mem_41__7__N_208), .Q(\mem[41] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i5 (.D(data[4]), .CK(mem_41__7__N_208), .Q(\mem[41] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i6 (.D(data[5]), .CK(mem_41__7__N_208), .Q(\mem[41] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i7 (.D(data[6]), .CK(mem_41__7__N_208), .Q(\mem[41] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i8 (.D(data[7]), .CK(mem_41__7__N_208), .Q(\mem[41] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i2 (.D(data[1]), .CK(mem_40__7__N_205), .Q(\mem[40] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i3 (.D(data[2]), .CK(mem_40__7__N_205), .Q(\mem[40] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i4 (.D(data[3]), .CK(mem_40__7__N_205), .Q(\mem[40] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i5 (.D(data[4]), .CK(mem_40__7__N_205), .Q(\mem[40] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i6 (.D(data[5]), .CK(mem_40__7__N_205), .Q(\mem[40] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i7 (.D(data[6]), .CK(mem_40__7__N_205), .Q(\mem[40] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i8 (.D(data[7]), .CK(mem_40__7__N_205), .Q(\mem[40] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i2 (.D(data[1]), .CK(mem_39__7__N_202), .Q(\mem[39] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i3 (.D(data[2]), .CK(mem_39__7__N_202), .Q(\mem[39] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i4 (.D(data[3]), .CK(mem_39__7__N_202), .Q(\mem[39] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i5 (.D(data[4]), .CK(mem_39__7__N_202), .Q(\mem[39] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i6 (.D(data[5]), .CK(mem_39__7__N_202), .Q(\mem[39] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i7 (.D(data[6]), .CK(mem_39__7__N_202), .Q(\mem[39] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i8 (.D(data[7]), .CK(mem_39__7__N_202), .Q(\mem[39] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i2 (.D(data[1]), .CK(mem_38__7__N_199), .Q(\mem[38] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i3 (.D(data[2]), .CK(mem_38__7__N_199), .Q(\mem[38] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i4 (.D(data[3]), .CK(mem_38__7__N_199), .Q(\mem[38] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i5 (.D(data[4]), .CK(mem_38__7__N_199), .Q(\mem[38] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i6 (.D(data[5]), .CK(mem_38__7__N_199), .Q(\mem[38] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i7 (.D(data[6]), .CK(mem_38__7__N_199), .Q(\mem[38] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i8 (.D(data[7]), .CK(mem_38__7__N_199), .Q(\mem[38] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i2 (.D(data[1]), .CK(mem_37__7__N_196), .Q(\mem[37] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i3 (.D(data[2]), .CK(mem_37__7__N_196), .Q(\mem[37] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i4 (.D(data[3]), .CK(mem_37__7__N_196), .Q(\mem[37] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i5 (.D(data[4]), .CK(mem_37__7__N_196), .Q(\mem[37] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i6 (.D(data[5]), .CK(mem_37__7__N_196), .Q(\mem[37] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i7 (.D(data[6]), .CK(mem_37__7__N_196), .Q(\mem[37] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i8 (.D(data[7]), .CK(mem_37__7__N_196), .Q(\mem[37] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i2 (.D(data[1]), .CK(mem_36__7__N_193), .Q(\mem[36] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i3 (.D(data[2]), .CK(mem_36__7__N_193), .Q(\mem[36] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i4 (.D(data[3]), .CK(mem_36__7__N_193), .Q(\mem[36] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i5 (.D(data[4]), .CK(mem_36__7__N_193), .Q(\mem[36] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i6 (.D(data[5]), .CK(mem_36__7__N_193), .Q(\mem[36] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i7 (.D(data[6]), .CK(mem_36__7__N_193), .Q(\mem[36] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i8 (.D(data[7]), .CK(mem_36__7__N_193), .Q(\mem[36] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i2 (.D(data[1]), .CK(mem_35__7__N_190), .Q(\mem[35] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i3 (.D(data[2]), .CK(mem_35__7__N_190), .Q(\mem[35] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i4 (.D(data[3]), .CK(mem_35__7__N_190), .Q(\mem[35] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i5 (.D(data[4]), .CK(mem_35__7__N_190), .Q(\mem[35] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i6 (.D(data[5]), .CK(mem_35__7__N_190), .Q(\mem[35] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i7 (.D(data[6]), .CK(mem_35__7__N_190), .Q(\mem[35] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i8 (.D(data[7]), .CK(mem_35__7__N_190), .Q(\mem[35] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i2 (.D(data[1]), .CK(mem_34__7__N_187), .Q(\mem[34] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i3 (.D(data[2]), .CK(mem_34__7__N_187), .Q(\mem[34] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i4 (.D(data[3]), .CK(mem_34__7__N_187), .Q(\mem[34] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i5 (.D(data[4]), .CK(mem_34__7__N_187), .Q(\mem[34] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i6 (.D(data[5]), .CK(mem_34__7__N_187), .Q(\mem[34] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i7 (.D(data[6]), .CK(mem_34__7__N_187), .Q(\mem[34] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i8 (.D(data[7]), .CK(mem_34__7__N_187), .Q(\mem[34] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i2 (.D(data[1]), .CK(mem_33__7__N_184), .Q(\mem[33] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i3 (.D(data[2]), .CK(mem_33__7__N_184), .Q(\mem[33] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i4 (.D(data[3]), .CK(mem_33__7__N_184), .Q(\mem[33] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i5 (.D(data[4]), .CK(mem_33__7__N_184), .Q(\mem[33] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i6 (.D(data[5]), .CK(mem_33__7__N_184), .Q(\mem[33] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i7 (.D(data[6]), .CK(mem_33__7__N_184), .Q(\mem[33] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i8 (.D(data[7]), .CK(mem_33__7__N_184), .Q(\mem[33] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i2 (.D(data[1]), .CK(mem_32__7__N_181), .Q(\mem[32] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i3 (.D(data[2]), .CK(mem_32__7__N_181), .Q(\mem[32] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i4 (.D(data[3]), .CK(mem_32__7__N_181), .Q(\mem[32] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i5 (.D(data[4]), .CK(mem_32__7__N_181), .Q(\mem[32] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i6 (.D(data[5]), .CK(mem_32__7__N_181), .Q(\mem[32] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i7 (.D(data[6]), .CK(mem_32__7__N_181), .Q(\mem[32] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i8 (.D(data[7]), .CK(mem_32__7__N_181), .Q(\mem[32] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i2 (.D(data[1]), .CK(mem_31__7__N_178), .Q(\mem[31] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i3 (.D(data[2]), .CK(mem_31__7__N_178), .Q(\mem[31] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i4 (.D(data[3]), .CK(mem_31__7__N_178), .Q(\mem[31] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i5 (.D(data[4]), .CK(mem_31__7__N_178), .Q(\mem[31] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i6 (.D(data[5]), .CK(mem_31__7__N_178), .Q(\mem[31] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i7 (.D(data[6]), .CK(mem_31__7__N_178), .Q(\mem[31] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i8 (.D(data[7]), .CK(mem_31__7__N_178), .Q(\mem[31] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i2 (.D(data[1]), .CK(mem_30__7__N_175), .Q(\mem[30] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i3 (.D(data[2]), .CK(mem_30__7__N_175), .Q(\mem[30] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i4 (.D(data[3]), .CK(mem_30__7__N_175), .Q(\mem[30] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i5 (.D(data[4]), .CK(mem_30__7__N_175), .Q(\mem[30] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i6 (.D(data[5]), .CK(mem_30__7__N_175), .Q(\mem[30] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i7 (.D(data[6]), .CK(mem_30__7__N_175), .Q(\mem[30] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i8 (.D(data[7]), .CK(mem_30__7__N_175), .Q(\mem[30] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i2 (.D(data[1]), .CK(mem_29__7__N_172), .Q(\mem[29] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i3 (.D(data[2]), .CK(mem_29__7__N_172), .Q(\mem[29] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i4 (.D(data[3]), .CK(mem_29__7__N_172), .Q(\mem[29] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i5 (.D(data[4]), .CK(mem_29__7__N_172), .Q(\mem[29] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i6 (.D(data[5]), .CK(mem_29__7__N_172), .Q(\mem[29] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i7 (.D(data[6]), .CK(mem_29__7__N_172), .Q(\mem[29] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i8 (.D(data[7]), .CK(mem_29__7__N_172), .Q(\mem[29] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i2 (.D(data[1]), .CK(mem_28__7__N_169), .Q(\mem[28] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i3 (.D(data[2]), .CK(mem_28__7__N_169), .Q(\mem[28] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i4 (.D(data[3]), .CK(mem_28__7__N_169), .Q(\mem[28] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i5 (.D(data[4]), .CK(mem_28__7__N_169), .Q(\mem[28] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i6 (.D(data[5]), .CK(mem_28__7__N_169), .Q(\mem[28] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i7 (.D(data[6]), .CK(mem_28__7__N_169), .Q(\mem[28] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i8 (.D(data[7]), .CK(mem_28__7__N_169), .Q(\mem[28] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i2 (.D(data[1]), .CK(mem_27__7__N_166), .Q(\mem[27] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i3 (.D(data[2]), .CK(mem_27__7__N_166), .Q(\mem[27] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i4 (.D(data[3]), .CK(mem_27__7__N_166), .Q(\mem[27] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i5 (.D(data[4]), .CK(mem_27__7__N_166), .Q(\mem[27] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i6 (.D(data[5]), .CK(mem_27__7__N_166), .Q(\mem[27] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i7 (.D(data[6]), .CK(mem_27__7__N_166), .Q(\mem[27] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i8 (.D(data[7]), .CK(mem_27__7__N_166), .Q(\mem[27] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i2 (.D(data[1]), .CK(mem_26__7__N_163), .Q(\mem[26] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i3 (.D(data[2]), .CK(mem_26__7__N_163), .Q(\mem[26] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i4 (.D(data[3]), .CK(mem_26__7__N_163), .Q(\mem[26] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i5 (.D(data[4]), .CK(mem_26__7__N_163), .Q(\mem[26] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i6 (.D(data[5]), .CK(mem_26__7__N_163), .Q(\mem[26] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i7 (.D(data[6]), .CK(mem_26__7__N_163), .Q(\mem[26] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i8 (.D(data[7]), .CK(mem_26__7__N_163), .Q(\mem[26] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i2 (.D(data[1]), .CK(mem_25__7__N_160), .Q(\mem[25] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i3 (.D(data[2]), .CK(mem_25__7__N_160), .Q(\mem[25] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i4 (.D(data[3]), .CK(mem_25__7__N_160), .Q(\mem[25] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i5 (.D(data[4]), .CK(mem_25__7__N_160), .Q(\mem[25] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i6 (.D(data[5]), .CK(mem_25__7__N_160), .Q(\mem[25] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i7 (.D(data[6]), .CK(mem_25__7__N_160), .Q(\mem[25] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i8 (.D(data[7]), .CK(mem_25__7__N_160), .Q(\mem[25] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i2 (.D(data[1]), .CK(mem_24__7__N_157), .Q(\mem[24] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i3 (.D(data[2]), .CK(mem_24__7__N_157), .Q(\mem[24] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i4 (.D(data[3]), .CK(mem_24__7__N_157), .Q(\mem[24] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i5 (.D(data[4]), .CK(mem_24__7__N_157), .Q(\mem[24] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i6 (.D(data[5]), .CK(mem_24__7__N_157), .Q(\mem[24] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i7 (.D(data[6]), .CK(mem_24__7__N_157), .Q(\mem[24] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i8 (.D(data[7]), .CK(mem_24__7__N_157), .Q(\mem[24] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i2 (.D(data[1]), .CK(mem_23__7__N_154), .Q(\mem[23] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i3 (.D(data[2]), .CK(mem_23__7__N_154), .Q(\mem[23] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i4 (.D(data[3]), .CK(mem_23__7__N_154), .Q(\mem[23] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i5 (.D(data[4]), .CK(mem_23__7__N_154), .Q(\mem[23] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i6 (.D(data[5]), .CK(mem_23__7__N_154), .Q(\mem[23] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i7 (.D(data[6]), .CK(mem_23__7__N_154), .Q(\mem[23] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i8 (.D(data[7]), .CK(mem_23__7__N_154), .Q(\mem[23] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i2 (.D(data[1]), .CK(mem_22__7__N_151), .Q(\mem[22] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i3 (.D(data[2]), .CK(mem_22__7__N_151), .Q(\mem[22] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i4 (.D(data[3]), .CK(mem_22__7__N_151), .Q(\mem[22] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i5 (.D(data[4]), .CK(mem_22__7__N_151), .Q(\mem[22] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i6 (.D(data[5]), .CK(mem_22__7__N_151), .Q(\mem[22] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i7 (.D(data[6]), .CK(mem_22__7__N_151), .Q(\mem[22] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i8 (.D(data[7]), .CK(mem_22__7__N_151), .Q(\mem[22] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i2 (.D(data[1]), .CK(mem_21__7__N_148), .Q(\mem[21] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i3 (.D(data[2]), .CK(mem_21__7__N_148), .Q(\mem[21] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i4 (.D(data[3]), .CK(mem_21__7__N_148), .Q(\mem[21] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i5 (.D(data[4]), .CK(mem_21__7__N_148), .Q(\mem[21] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i6 (.D(data[5]), .CK(mem_21__7__N_148), .Q(\mem[21] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i7 (.D(data[6]), .CK(mem_21__7__N_148), .Q(\mem[21] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i8 (.D(data[7]), .CK(mem_21__7__N_148), .Q(\mem[21] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i8.GSR = "DISABLED";
    LUT4 i1459_3_lut (.A(\mem[28] [7]), .B(\mem[29] [7]), .C(address[0]), 
         .Z(n1529)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1459_3_lut.init = 16'hcaca;
    PFUMX i1528 (.BLUT(n1587), .ALUT(n1588), .C0(address[1]), .Z(n1598));
    PFUMX i1403 (.BLUT(n1461), .ALUT(n1462), .C0(address[1]), .Z(n1473));
    PFUMX i1368 (.BLUT(n1422), .ALUT(n1423), .C0(address[1]), .Z(n1438));
    PFUMX i1404 (.BLUT(n1463), .ALUT(n1464), .C0(address[1]), .Z(n1474));
    LUT4 i1458_3_lut (.A(\mem[26] [7]), .B(\mem[27] [7]), .C(address[0]), 
         .Z(n1528)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1458_3_lut.init = 16'hcaca;
    PFUMX i1400 (.BLUT(n1455), .ALUT(n1456), .C0(address[1]), .Z(n1470));
    LUT4 i1582_3_lut (.A(\mem[58] [6]), .B(\mem[59] [6]), .C(address[0]), 
         .Z(n1652)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1582_3_lut.init = 16'hcaca;
    PFUMX i1466 (.BLUT(n1525), .ALUT(n1526), .C0(address[1]), .Z(n1536));
    PFUMX i1560 (.BLUT(n1620), .ALUT(n1621), .C0(address[1]), .Z(n1630));
    PFUMX i1561 (.BLUT(n1622), .ALUT(n1623), .C0(address[1]), .Z(n1631));
    PFUMX i1405 (.BLUT(n1465), .ALUT(n1466), .C0(address[1]), .Z(n1475));
    LUT4 i1581_3_lut (.A(\mem[56] [6]), .B(\mem[57] [6]), .C(address[0]), 
         .Z(n1651)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1581_3_lut.init = 16'hcaca;
    PFUMX i1467 (.BLUT(n1527), .ALUT(n1528), .C0(address[1]), .Z(n1537));
    LUT4 i1429_3_lut (.A(\mem[30] [0]), .B(\mem[31] [0]), .C(address[0]), 
         .Z(n1499)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1429_3_lut.init = 16'hcaca;
    PFUMX i1652 (.BLUT(n1711), .ALUT(n1712), .C0(address[1]), .Z(n1722));
    LUT4 i1428_3_lut (.A(\mem[28] [0]), .B(\mem[29] [0]), .C(address[0]), 
         .Z(n1498)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1428_3_lut.init = 16'hcaca;
    LUT4 i1427_3_lut (.A(\mem[26] [0]), .B(\mem[27] [0]), .C(address[0]), 
         .Z(n1497)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1427_3_lut.init = 16'hcaca;
    LUT4 i1426_3_lut (.A(\mem[24] [0]), .B(\mem[25] [0]), .C(address[0]), 
         .Z(n1496)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1426_3_lut.init = 16'hcaca;
    PFUMX i1401 (.BLUT(n1457), .ALUT(n1458), .C0(address[1]), .Z(n1471));
    PFUMX i1369 (.BLUT(n1424), .ALUT(n1425), .C0(address[1]), .Z(n1439));
    PFUMX i1406 (.BLUT(n1467), .ALUT(n1468), .C0(address[1]), .Z(n1476));
    LUT4 i1580_3_lut (.A(\mem[54] [6]), .B(\mem[55] [6]), .C(address[0]), 
         .Z(n1650)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1580_3_lut.init = 16'hcaca;
    LUT4 i1579_3_lut (.A(\mem[52] [6]), .B(\mem[53] [6]), .C(address[0]), 
         .Z(n1649)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1579_3_lut.init = 16'hcaca;
    LUT4 i1425_3_lut (.A(\mem[22] [0]), .B(\mem[23] [0]), .C(address[0]), 
         .Z(n1495)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1425_3_lut.init = 16'hcaca;
    PFUMX i1653 (.BLUT(n1713), .ALUT(n1714), .C0(address[1]), .Z(n1723));
    LUT4 i1424_3_lut (.A(\mem[20] [0]), .B(\mem[21] [0]), .C(address[0]), 
         .Z(n1494)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1424_3_lut.init = 16'hcaca;
    PFUMX i1654 (.BLUT(n1715), .ALUT(n1716), .C0(address[1]), .Z(n1724));
    LUT4 i1423_3_lut (.A(\mem[18] [0]), .B(\mem[19] [0]), .C(address[0]), 
         .Z(n1493)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1423_3_lut.init = 16'hcaca;
    LUT4 i1422_3_lut (.A(\mem[16] [0]), .B(\mem[17] [0]), .C(address[0]), 
         .Z(n1492)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1422_3_lut.init = 16'hcaca;
    PFUMX i1244 (.BLUT(n1298), .ALUT(n1299), .C0(address[1]), .Z(n1314));
    LUT4 Select_348_i3_4_lut (.A(data_7__N_66[0]), .B(akku_o_c_0), .C(data_7__N_79), 
         .D(n1891), .Z(data[0])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_348_i3_4_lut.init = 16'ha0ec;
    LUT4 i1578_3_lut (.A(\mem[50] [6]), .B(\mem[51] [6]), .C(address[0]), 
         .Z(n1648)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1578_3_lut.init = 16'hcaca;
    PFUMX i1251 (.BLUT(n1312), .ALUT(n1313), .C0(address[1]), .Z(n1321));
    LUT4 i1577_3_lut (.A(\mem[48] [6]), .B(\mem[49] [6]), .C(address[0]), 
         .Z(n1647)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1577_3_lut.init = 16'hcaca;
    LUT4 i1421_3_lut (.A(\mem[14] [0]), .B(\mem[15] [0]), .C(address[0]), 
         .Z(n1491)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1421_3_lut.init = 16'hcaca;
    LUT4 i1420_3_lut (.A(\mem[12] [0]), .B(\mem[13] [0]), .C(address[0]), 
         .Z(n1490)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1420_3_lut.init = 16'hcaca;
    PFUMX i1245 (.BLUT(n1300), .ALUT(n1301), .C0(address[1]), .Z(n1315));
    PFUMX i1530 (.BLUT(n1591), .ALUT(n1592), .C0(address[1]), .Z(n1600));
    LUT4 i1475_3_lut (.A(n1543), .B(n1544), .C(address[4]), .Z(n1545)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1475_3_lut.init = 16'hcaca;
    LUT4 i1506_3_lut (.A(n1574), .B(n1575), .C(address[4]), .Z(n1576)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1506_3_lut.init = 16'hcaca;
    LUT4 i1444_3_lut (.A(n1512), .B(n1513), .C(address[4]), .Z(n1514)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1444_3_lut.init = 16'hcaca;
    LUT4 i1537_3_lut (.A(n1605), .B(n1606), .C(address[4]), .Z(n1607)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1537_3_lut.init = 16'hcaca;
    LUT4 i1413_3_lut (.A(n1481), .B(n1482), .C(address[4]), .Z(n1483)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1413_3_lut.init = 16'hcaca;
    LUT4 i1568_3_lut (.A(n1636), .B(n1637), .C(address[4]), .Z(n1638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1568_3_lut.init = 16'hcaca;
    LUT4 i1382_3_lut (.A(n1450), .B(n1451), .C(address[4]), .Z(n1452)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1382_3_lut.init = 16'hcaca;
    LUT4 i1599_3_lut (.A(n1667), .B(n1668), .C(address[4]), .Z(n1669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1599_3_lut.init = 16'hcaca;
    LUT4 i1351_3_lut (.A(n1419), .B(n1420), .C(address[4]), .Z(n1421)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1351_3_lut.init = 16'hcaca;
    LUT4 i1630_3_lut (.A(n1698), .B(n1699), .C(address[4]), .Z(n1700)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1630_3_lut.init = 16'hcaca;
    LUT4 i1320_3_lut (.A(n1388), .B(n1389), .C(address[4]), .Z(n1390)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1320_3_lut.init = 16'hcaca;
    LUT4 i1419_3_lut (.A(\mem[10] [0]), .B(\mem[11] [0]), .C(address[0]), 
         .Z(n1489)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1419_3_lut.init = 16'hcaca;
    PFUMX i1246 (.BLUT(n1302), .ALUT(n1303), .C0(address[1]), .Z(n1316));
    LUT4 i1661_3_lut (.A(n1729), .B(n1730), .C(address[4]), .Z(n1731)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1661_3_lut.init = 16'hcaca;
    LUT4 i1289_3_lut (.A(n1357), .B(n1358), .C(address[4]), .Z(n1359)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1289_3_lut.init = 16'hcaca;
    LUT4 i1692_3_lut (.A(n1760), .B(n1761), .C(address[4]), .Z(n1762)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1692_3_lut.init = 16'hcaca;
    LUT4 i1258_3_lut (.A(n1326), .B(n1327), .C(address[4]), .Z(n1328)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1258_3_lut.init = 16'hcaca;
    LUT4 i1723_3_lut (.A(n1791), .B(n1792), .C(address[4]), .Z(n1793)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1723_3_lut.init = 16'hcaca;
    LUT4 i1259_3_lut (.A(\mem[0] [5]), .B(\mem[1] [5]), .C(address[0]), 
         .Z(n1329)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1259_3_lut.init = 16'hcaca;
    LUT4 i1260_3_lut (.A(\mem[2] [5]), .B(\mem[3] [5]), .C(address[0]), 
         .Z(n1330)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1260_3_lut.init = 16'hcaca;
    LUT4 i1261_3_lut (.A(\mem[4] [5]), .B(\mem[5] [5]), .C(address[0]), 
         .Z(n1331)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1261_3_lut.init = 16'hcaca;
    LUT4 i1262_3_lut (.A(\mem[6] [5]), .B(\mem[7] [5]), .C(address[0]), 
         .Z(n1332)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1262_3_lut.init = 16'hcaca;
    LUT4 i1418_3_lut (.A(\mem[8] [0]), .B(\mem[9] [0]), .C(address[0]), 
         .Z(n1488)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1418_3_lut.init = 16'hcaca;
    LUT4 i1263_3_lut (.A(\mem[8] [5]), .B(\mem[9] [5]), .C(address[0]), 
         .Z(n1333)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1263_3_lut.init = 16'hcaca;
    LUT4 i1264_3_lut (.A(\mem[10] [5]), .B(\mem[11] [5]), .C(address[0]), 
         .Z(n1334)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1264_3_lut.init = 16'hcaca;
    LUT4 i1265_3_lut (.A(\mem[12] [5]), .B(\mem[13] [5]), .C(address[0]), 
         .Z(n1335)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1265_3_lut.init = 16'hcaca;
    LUT4 i1266_3_lut (.A(\mem[14] [5]), .B(\mem[15] [5]), .C(address[0]), 
         .Z(n1336)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1266_3_lut.init = 16'hcaca;
    LUT4 i1267_3_lut (.A(\mem[16] [5]), .B(\mem[17] [5]), .C(address[0]), 
         .Z(n1337)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1267_3_lut.init = 16'hcaca;
    LUT4 i1268_3_lut (.A(\mem[18] [5]), .B(\mem[19] [5]), .C(address[0]), 
         .Z(n1338)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1268_3_lut.init = 16'hcaca;
    LUT4 i1269_3_lut (.A(\mem[20] [5]), .B(\mem[21] [5]), .C(address[0]), 
         .Z(n1339)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1269_3_lut.init = 16'hcaca;
    LUT4 i1270_3_lut (.A(\mem[22] [5]), .B(\mem[23] [5]), .C(address[0]), 
         .Z(n1340)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1270_3_lut.init = 16'hcaca;
    LUT4 i1271_3_lut (.A(\mem[24] [5]), .B(\mem[25] [5]), .C(address[0]), 
         .Z(n1341)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1271_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_69 (.A(address[4]), .B(address[3]), .C(address[5]), 
         .Z(n684)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_adj_69.init = 16'hf7f7;
    LUT4 i1272_3_lut (.A(\mem[26] [5]), .B(\mem[27] [5]), .C(address[0]), 
         .Z(n1342)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1272_3_lut.init = 16'hcaca;
    LUT4 i1273_3_lut (.A(\mem[28] [5]), .B(\mem[29] [5]), .C(address[0]), 
         .Z(n1343)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1273_3_lut.init = 16'hcaca;
    LUT4 i1274_3_lut (.A(\mem[30] [5]), .B(\mem[31] [5]), .C(address[0]), 
         .Z(n1344)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1274_3_lut.init = 16'hcaca;
    LUT4 i1666_3_lut (.A(\mem[40] [5]), .B(\mem[41] [5]), .C(address[0]), 
         .Z(n1736)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1666_3_lut.init = 16'hcaca;
    LUT4 i1667_3_lut (.A(\mem[42] [5]), .B(\mem[43] [5]), .C(address[0]), 
         .Z(n1737)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1667_3_lut.init = 16'hcaca;
    LUT4 i1600_3_lut (.A(\mem[32] [3]), .B(\mem[33] [3]), .C(address[0]), 
         .Z(n1670)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1600_3_lut.init = 16'hcaca;
    LUT4 i1601_3_lut (.A(\mem[34] [3]), .B(\mem[35] [3]), .C(address[0]), 
         .Z(n1671)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1601_3_lut.init = 16'hcaca;
    LUT4 i1602_3_lut (.A(\mem[36] [3]), .B(\mem[37] [3]), .C(address[0]), 
         .Z(n1672)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1602_3_lut.init = 16'hcaca;
    LUT4 i1603_3_lut (.A(\mem[38] [3]), .B(\mem[39] [3]), .C(address[0]), 
         .Z(n1673)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1603_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_70 (.A(address[4]), .B(address[3]), .C(address[5]), 
         .Z(n1272)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_70.init = 16'h8080;
    PFUMX i1247 (.BLUT(n1304), .ALUT(n1305), .C0(address[1]), .Z(n1317));
    LUT4 i1476_3_lut (.A(\mem[32] [7]), .B(\mem[33] [7]), .C(address[0]), 
         .Z(n1546)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1476_3_lut.init = 16'hcaca;
    LUT4 i1477_3_lut (.A(\mem[34] [7]), .B(\mem[35] [7]), .C(address[0]), 
         .Z(n1547)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1477_3_lut.init = 16'hcaca;
    LUT4 i1604_3_lut (.A(\mem[40] [3]), .B(\mem[41] [3]), .C(address[0]), 
         .Z(n1674)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1604_3_lut.init = 16'hcaca;
    LUT4 i1605_3_lut (.A(\mem[42] [3]), .B(\mem[43] [3]), .C(address[0]), 
         .Z(n1675)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1605_3_lut.init = 16'hcaca;
    LUT4 i1668_3_lut (.A(\mem[44] [5]), .B(\mem[45] [5]), .C(address[0]), 
         .Z(n1738)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1668_3_lut.init = 16'hcaca;
    LUT4 i1669_3_lut (.A(\mem[46] [5]), .B(\mem[47] [5]), .C(address[0]), 
         .Z(n1739)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1669_3_lut.init = 16'hcaca;
    LUT4 i1701_3_lut (.A(\mem[48] [1]), .B(\mem[49] [1]), .C(address[0]), 
         .Z(n1771)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1701_3_lut.init = 16'hcaca;
    LUT4 i1702_3_lut (.A(\mem[50] [1]), .B(\mem[51] [1]), .C(address[0]), 
         .Z(n1772)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1702_3_lut.init = 16'hcaca;
    LUT4 i1478_3_lut (.A(\mem[36] [7]), .B(\mem[37] [7]), .C(address[0]), 
         .Z(n1548)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1478_3_lut.init = 16'hcaca;
    PFUMX i1679 (.BLUT(n1734), .ALUT(n1735), .C0(address[1]), .Z(n1749));
    LUT4 i1479_3_lut (.A(\mem[38] [7]), .B(\mem[39] [7]), .C(address[0]), 
         .Z(n1549)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1479_3_lut.init = 16'hcaca;
    LUT4 i1480_3_lut (.A(\mem[40] [7]), .B(\mem[41] [7]), .C(address[0]), 
         .Z(n1550)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1480_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut (.A(n1896), .B(n1890), .C(address[1]), .D(n1283), 
         .Z(mem_55__7__N_250)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0080;
    LUT4 i1481_3_lut (.A(\mem[42] [7]), .B(\mem[43] [7]), .C(address[0]), 
         .Z(n1551)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1481_3_lut.init = 16'hcaca;
    LUT4 i1606_3_lut (.A(\mem[44] [3]), .B(\mem[45] [3]), .C(address[0]), 
         .Z(n1676)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1606_3_lut.init = 16'hcaca;
    LUT4 i1607_3_lut (.A(\mem[46] [3]), .B(\mem[47] [3]), .C(address[0]), 
         .Z(n1677)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1607_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_71 (.A(n1896), .B(n1890), .C(address[1]), 
         .D(n1260), .Z(mem_47__7__N_226)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_71.init = 16'h0080;
    LUT4 i1_2_lut_4_lut_adj_72 (.A(n1896), .B(n1890), .C(address[1]), 
         .D(n1284), .Z(mem_39__7__N_202)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_72.init = 16'h0080;
    LUT4 i1482_3_lut (.A(\mem[44] [7]), .B(\mem[45] [7]), .C(address[0]), 
         .Z(n1552)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1482_3_lut.init = 16'hcaca;
    LUT4 i1483_3_lut (.A(\mem[46] [7]), .B(\mem[47] [7]), .C(address[0]), 
         .Z(n1553)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1483_3_lut.init = 16'hcaca;
    LUT4 i1484_3_lut (.A(\mem[48] [7]), .B(\mem[49] [7]), .C(address[0]), 
         .Z(n1554)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1484_3_lut.init = 16'hcaca;
    LUT4 i1485_3_lut (.A(\mem[50] [7]), .B(\mem[51] [7]), .C(address[0]), 
         .Z(n1555)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1485_3_lut.init = 16'hcaca;
    LUT4 i1608_3_lut (.A(\mem[48] [3]), .B(\mem[49] [3]), .C(address[0]), 
         .Z(n1678)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1608_3_lut.init = 16'hcaca;
    LUT4 i1609_3_lut (.A(\mem[50] [3]), .B(\mem[51] [3]), .C(address[0]), 
         .Z(n1679)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1609_3_lut.init = 16'hcaca;
    LUT4 i1670_3_lut (.A(\mem[48] [5]), .B(\mem[49] [5]), .C(address[0]), 
         .Z(n1740)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1670_3_lut.init = 16'hcaca;
    LUT4 i1671_3_lut (.A(\mem[50] [5]), .B(\mem[51] [5]), .C(address[0]), 
         .Z(n1741)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1671_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_73 (.A(n1896), .B(n1890), .C(address[1]), 
         .D(n684), .Z(mem_31__7__N_178)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_73.init = 16'h0080;
    PFUMX i1370 (.BLUT(n1426), .ALUT(n1427), .C0(address[1]), .Z(n1440));
    LUT4 i1290_3_lut (.A(\mem[0] [4]), .B(\mem[1] [4]), .C(address[0]), 
         .Z(n1360)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1290_3_lut.init = 16'hcaca;
    LUT4 i1291_3_lut (.A(\mem[2] [4]), .B(\mem[3] [4]), .C(address[0]), 
         .Z(n1361)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1291_3_lut.init = 16'hcaca;
    LUT4 i1486_3_lut (.A(\mem[52] [7]), .B(\mem[53] [7]), .C(address[0]), 
         .Z(n1556)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1486_3_lut.init = 16'hcaca;
    LUT4 i1487_3_lut (.A(\mem[54] [7]), .B(\mem[55] [7]), .C(address[0]), 
         .Z(n1557)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1487_3_lut.init = 16'hcaca;
    LUT4 i1292_3_lut (.A(\mem[4] [4]), .B(\mem[5] [4]), .C(address[0]), 
         .Z(n1362)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1292_3_lut.init = 16'hcaca;
    LUT4 i1293_3_lut (.A(\mem[6] [4]), .B(\mem[7] [4]), .C(address[0]), 
         .Z(n1363)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1293_3_lut.init = 16'hcaca;
    LUT4 i1488_3_lut (.A(\mem[56] [7]), .B(\mem[57] [7]), .C(address[0]), 
         .Z(n1558)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1488_3_lut.init = 16'hcaca;
    LUT4 i1489_3_lut (.A(\mem[58] [7]), .B(\mem[59] [7]), .C(address[0]), 
         .Z(n1559)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1489_3_lut.init = 16'hcaca;
    LUT4 i1610_3_lut (.A(\mem[52] [3]), .B(\mem[53] [3]), .C(address[0]), 
         .Z(n1680)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1610_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_74 (.A(n1896), .B(n1890), .C(address[1]), 
         .D(n1261), .Z(mem_23__7__N_154)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_74.init = 16'h0080;
    LUT4 i1611_3_lut (.A(\mem[54] [3]), .B(\mem[55] [3]), .C(address[0]), 
         .Z(n1681)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1611_3_lut.init = 16'hcaca;
    LUT4 i1294_3_lut (.A(\mem[8] [4]), .B(\mem[9] [4]), .C(address[0]), 
         .Z(n1364)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1294_3_lut.init = 16'hcaca;
    LUT4 i1295_3_lut (.A(\mem[10] [4]), .B(\mem[11] [4]), .C(address[0]), 
         .Z(n1365)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1295_3_lut.init = 16'hcaca;
    LUT4 i1296_3_lut (.A(\mem[12] [4]), .B(\mem[13] [4]), .C(address[0]), 
         .Z(n1366)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1296_3_lut.init = 16'hcaca;
    LUT4 i1297_3_lut (.A(\mem[14] [4]), .B(\mem[15] [4]), .C(address[0]), 
         .Z(n1367)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1297_3_lut.init = 16'hcaca;
    LUT4 i1490_3_lut (.A(\mem[60] [7]), .B(\mem[61] [7]), .C(address[0]), 
         .Z(n1560)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1490_3_lut.init = 16'hcaca;
    LUT4 i1491_3_lut (.A(\mem[62] [7]), .B(\mem[63] [7]), .C(address[0]), 
         .Z(n1561)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1491_3_lut.init = 16'hcaca;
    LUT4 i1612_3_lut (.A(\mem[56] [3]), .B(\mem[57] [3]), .C(address[0]), 
         .Z(n1682)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1612_3_lut.init = 16'hcaca;
    LUT4 i1613_3_lut (.A(\mem[58] [3]), .B(\mem[59] [3]), .C(address[0]), 
         .Z(n1683)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1613_3_lut.init = 16'hcaca;
    LUT4 i1672_3_lut (.A(\mem[52] [5]), .B(\mem[53] [5]), .C(address[0]), 
         .Z(n1742)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1672_3_lut.init = 16'hcaca;
    LUT4 i1673_3_lut (.A(\mem[54] [5]), .B(\mem[55] [5]), .C(address[0]), 
         .Z(n1743)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1673_3_lut.init = 16'hcaca;
    LUT4 i1298_3_lut (.A(\mem[16] [4]), .B(\mem[17] [4]), .C(address[0]), 
         .Z(n1368)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1298_3_lut.init = 16'hcaca;
    LUT4 i1299_3_lut (.A(\mem[18] [4]), .B(\mem[19] [4]), .C(address[0]), 
         .Z(n1369)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1299_3_lut.init = 16'hcaca;
    LUT4 i1300_3_lut (.A(\mem[20] [4]), .B(\mem[21] [4]), .C(address[0]), 
         .Z(n1370)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1300_3_lut.init = 16'hcaca;
    LUT4 i1301_3_lut (.A(\mem[22] [4]), .B(\mem[23] [4]), .C(address[0]), 
         .Z(n1371)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1301_3_lut.init = 16'hcaca;
    LUT4 i1302_3_lut (.A(\mem[24] [4]), .B(\mem[25] [4]), .C(address[0]), 
         .Z(n1372)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1302_3_lut.init = 16'hcaca;
    LUT4 i1303_3_lut (.A(\mem[26] [4]), .B(\mem[27] [4]), .C(address[0]), 
         .Z(n1373)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1303_3_lut.init = 16'hcaca;
    LUT4 i1304_3_lut (.A(\mem[28] [4]), .B(\mem[29] [4]), .C(address[0]), 
         .Z(n1374)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1304_3_lut.init = 16'hcaca;
    PFUMX i1371 (.BLUT(n1428), .ALUT(n1429), .C0(address[1]), .Z(n1441));
    LUT4 i1305_3_lut (.A(\mem[30] [4]), .B(\mem[31] [4]), .C(address[0]), 
         .Z(n1375)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1305_3_lut.init = 16'hcaca;
    LUT4 i1614_3_lut (.A(\mem[60] [3]), .B(\mem[61] [3]), .C(address[0]), 
         .Z(n1684)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1614_3_lut.init = 16'hcaca;
    LUT4 i1615_3_lut (.A(\mem[62] [3]), .B(\mem[63] [3]), .C(address[0]), 
         .Z(n1685)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1615_3_lut.init = 16'hcaca;
    LUT4 i1674_3_lut (.A(\mem[56] [5]), .B(\mem[57] [5]), .C(address[0]), 
         .Z(n1744)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1674_3_lut.init = 16'hcaca;
    LUT4 i1675_3_lut (.A(\mem[58] [5]), .B(\mem[59] [5]), .C(address[0]), 
         .Z(n1745)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1675_3_lut.init = 16'hcaca;
    LUT4 i1703_3_lut (.A(\mem[52] [1]), .B(\mem[53] [1]), .C(address[0]), 
         .Z(n1773)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1703_3_lut.init = 16'hcaca;
    LUT4 i1704_3_lut (.A(\mem[54] [1]), .B(\mem[55] [1]), .C(address[0]), 
         .Z(n1774)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1704_3_lut.init = 16'hcaca;
    LUT4 i1236_3_lut (.A(\mem[16] [1]), .B(\mem[17] [1]), .C(address[0]), 
         .Z(n1306)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1236_3_lut.init = 16'hcaca;
    LUT4 i1237_3_lut (.A(\mem[18] [1]), .B(\mem[19] [1]), .C(address[0]), 
         .Z(n1307)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1237_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut (.A(address[5]), .B(address[3]), .C(address[4]), .Z(n1260)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i2_3_lut.init = 16'hf7f7;
    LUT4 i1676_3_lut (.A(\mem[60] [5]), .B(\mem[61] [5]), .C(address[0]), 
         .Z(n1746)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1676_3_lut.init = 16'hcaca;
    LUT4 i1677_3_lut (.A(\mem[62] [5]), .B(\mem[63] [5]), .C(address[0]), 
         .Z(n1747)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1677_3_lut.init = 16'hcaca;
    LUT4 i1705_3_lut (.A(\mem[56] [1]), .B(\mem[57] [1]), .C(address[0]), 
         .Z(n1775)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1705_3_lut.init = 16'hcaca;
    LUT4 i1706_3_lut (.A(\mem[58] [1]), .B(\mem[59] [1]), .C(address[0]), 
         .Z(n1776)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1706_3_lut.init = 16'hcaca;
    LUT4 i1707_3_lut (.A(\mem[60] [1]), .B(\mem[61] [1]), .C(address[0]), 
         .Z(n1777)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1707_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_75 (.A(n1896), .B(n1890), .C(address[1]), 
         .D(n1272), .Z(mem_63__7__N_274)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_75.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_adj_76 (.A(address[0]), .B(address[1]), .C(address[2]), 
         .Z(n1295)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_adj_76.init = 16'hfefe;
    LUT4 i889_2_lut_rep_79 (.A(address[0]), .B(address[2]), .Z(n1896)) /* synthesis lut_function=(A (B)) */ ;
    defparam i889_2_lut_rep_79.init = 16'h8888;
    LUT4 i1569_3_lut (.A(\mem[32] [6]), .B(\mem[33] [6]), .C(address[0]), 
         .Z(n1639)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1569_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_77 (.A(n1896), .B(n1890), .C(address[1]), 
         .D(n1290), .Z(mem_15__7__N_130)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_77.init = 16'h0080;
    PFUMX i1372 (.BLUT(n1430), .ALUT(n1431), .C0(address[1]), .Z(n1442));
    LUT4 i1_2_lut_3_lut_adj_78 (.A(address[0]), .B(address[2]), .C(address[1]), 
         .Z(n681)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_adj_78.init = 16'hf7f7;
    LUT4 i1_2_lut_4_lut_adj_79 (.A(n1896), .B(n1890), .C(address[1]), 
         .D(n1289), .Z(mem_7__7__N_106)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_79.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_adj_80 (.A(address[0]), .B(address[1]), .C(address[2]), 
         .Z(n1287)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_adj_80.init = 16'hbfbf;
    LUT4 i1_2_lut_3_lut_adj_81 (.A(address[0]), .B(address[1]), .C(address[2]), 
         .Z(n1286)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_adj_81.init = 16'hfbfb;
    LUT4 i1576_3_lut (.A(\mem[46] [6]), .B(\mem[47] [6]), .C(address[0]), 
         .Z(n1646)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1576_3_lut.init = 16'hcaca;
    PFUMX i1373 (.BLUT(n1432), .ALUT(n1433), .C0(address[1]), .Z(n1443));
    LUT4 i1367_3_lut (.A(\mem[30] [6]), .B(\mem[31] [6]), .C(address[0]), 
         .Z(n1437)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1367_3_lut.init = 16'hcaca;
    LUT4 i1575_3_lut (.A(\mem[44] [6]), .B(\mem[45] [6]), .C(address[0]), 
         .Z(n1645)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1575_3_lut.init = 16'hcaca;
    LUT4 i1366_3_lut (.A(\mem[28] [6]), .B(\mem[29] [6]), .C(address[0]), 
         .Z(n1436)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1366_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_adj_82 (.A(address[4]), .B(address[5]), .C(address[3]), 
         .Z(n1261)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i2_3_lut_adj_82.init = 16'hfdfd;
    LUT4 i1417_3_lut (.A(\mem[6] [0]), .B(\mem[7] [0]), .C(address[0]), 
         .Z(n1487)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1417_3_lut.init = 16'hcaca;
    LUT4 i1416_3_lut (.A(\mem[4] [0]), .B(\mem[5] [0]), .C(address[0]), 
         .Z(n1486)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1416_3_lut.init = 16'hcaca;
    PFUMX i1374 (.BLUT(n1434), .ALUT(n1435), .C0(address[1]), .Z(n1444));
    LUT4 i1365_3_lut (.A(\mem[26] [6]), .B(\mem[27] [6]), .C(address[0]), 
         .Z(n1435)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1365_3_lut.init = 16'hcaca;
    LUT4 i1364_3_lut (.A(\mem[24] [6]), .B(\mem[25] [6]), .C(address[0]), 
         .Z(n1434)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1364_3_lut.init = 16'hcaca;
    LUT4 i1415_3_lut (.A(\mem[2] [0]), .B(\mem[3] [0]), .C(address[0]), 
         .Z(n1485)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1415_3_lut.init = 16'hcaca;
    LUT4 i1363_3_lut (.A(\mem[22] [6]), .B(\mem[23] [6]), .C(address[0]), 
         .Z(n1433)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1363_3_lut.init = 16'hcaca;
    LUT4 i1362_3_lut (.A(\mem[20] [6]), .B(\mem[21] [6]), .C(address[0]), 
         .Z(n1432)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1362_3_lut.init = 16'hcaca;
    LUT4 i1518_3_lut (.A(\mem[54] [0]), .B(\mem[55] [0]), .C(address[0]), 
         .Z(n1588)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1518_3_lut.init = 16'hcaca;
    PFUMX i1375 (.BLUT(n1436), .ALUT(n1437), .C0(address[1]), .Z(n1445));
    LUT4 Select_347_i3_4_lut (.A(data_7__N_66[1]), .B(akku_o_c_1), .C(data_7__N_79), 
         .D(n1891), .Z(data[1])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_347_i3_4_lut.init = 16'ha0ec;
    LUT4 Select_346_i3_4_lut (.A(data_7__N_66[2]), .B(akku_o_c_2), .C(data_7__N_79), 
         .D(n1891), .Z(data[2])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_346_i3_4_lut.init = 16'ha0ec;
    PFUMX i1529 (.BLUT(n1589), .ALUT(n1590), .C0(address[1]), .Z(n1599));
    LUT4 i1414_3_lut (.A(\mem[0] [0]), .B(\mem[1] [0]), .C(address[0]), 
         .Z(n1484)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1414_3_lut.init = 16'hcaca;
    LUT4 Select_345_i3_4_lut (.A(data_7__N_66[3]), .B(akku_o_c_3), .C(data_7__N_79), 
         .D(n1891), .Z(data[3])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_345_i3_4_lut.init = 16'ha0ec;
    LUT4 Select_344_i3_4_lut (.A(data_7__N_66[4]), .B(akku_o_c_4), .C(data_7__N_79), 
         .D(n1891), .Z(data[4])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_344_i3_4_lut.init = 16'ha0ec;
    LUT4 Select_343_i3_4_lut (.A(data_7__N_66[5]), .B(akku_o_c_5), .C(data_7__N_79), 
         .D(n1891), .Z(data[5])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_343_i3_4_lut.init = 16'ha0ec;
    LUT4 Select_342_i3_4_lut (.A(data_7__N_66[6]), .B(akku_o_c_6), .C(data_7__N_79), 
         .D(n1891), .Z(data[6])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_342_i3_4_lut.init = 16'ha0ec;
    LUT4 Select_341_i3_4_lut (.A(data_7__N_66[7]), .B(akku_o_c_7), .C(data_7__N_79), 
         .D(n1891), .Z(data[7])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_341_i3_4_lut.init = 16'ha0ec;
    LUT4 i1361_3_lut (.A(\mem[18] [6]), .B(\mem[19] [6]), .C(address[0]), 
         .Z(n1431)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1361_3_lut.init = 16'hcaca;
    LUT4 i1519_3_lut (.A(\mem[56] [0]), .B(\mem[57] [0]), .C(address[0]), 
         .Z(n1589)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1519_3_lut.init = 16'hcaca;
    LUT4 i1665_3_lut (.A(\mem[38] [5]), .B(\mem[39] [5]), .C(address[0]), 
         .Z(n1735)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1665_3_lut.init = 16'hcaca;
    PFUMX i1585 (.BLUT(n1639), .ALUT(n1640), .C0(address[1]), .Z(n1655));
    LUT4 i341_1_lut (.A(address[0]), .Z(\pc_5__N_30[0] )) /* synthesis lut_function=(!(A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i341_1_lut.init = 16'h5555;
    LUT4 i1664_3_lut (.A(\mem[36] [5]), .B(\mem[37] [5]), .C(address[0]), 
         .Z(n1734)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1664_3_lut.init = 16'hcaca;
    LUT4 i1360_3_lut (.A(\mem[16] [6]), .B(\mem[17] [6]), .C(address[0]), 
         .Z(n1430)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1360_3_lut.init = 16'hcaca;
    PFUMX i1402 (.BLUT(n1459), .ALUT(n1460), .C0(address[1]), .Z(n1472));
    PFUMX i1586 (.BLUT(n1641), .ALUT(n1642), .C0(address[1]), .Z(n1656));
    PFUMX i1587 (.BLUT(n1643), .ALUT(n1644), .C0(address[1]), .Z(n1657));
    PFUMX i1430 (.BLUT(n1484), .ALUT(n1485), .C0(address[1]), .Z(n1500));
    PFUMX i1431 (.BLUT(n1486), .ALUT(n1487), .C0(address[1]), .Z(n1501));
    PFUMX i1588 (.BLUT(n1645), .ALUT(n1646), .C0(address[1]), .Z(n1658));
    LUT4 i1359_3_lut (.A(\mem[14] [6]), .B(\mem[15] [6]), .C(address[0]), 
         .Z(n1429)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1359_3_lut.init = 16'hcaca;
    PFUMX i1249 (.BLUT(n1308), .ALUT(n1309), .C0(address[1]), .Z(n1319));
    LUT4 i1358_3_lut (.A(\mem[12] [6]), .B(\mem[13] [6]), .C(address[0]), 
         .Z(n1428)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1358_3_lut.init = 16'hcaca;
    LUT4 i1357_3_lut (.A(\mem[10] [6]), .B(\mem[11] [6]), .C(address[0]), 
         .Z(n1427)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1357_3_lut.init = 16'hcaca;
    LUT4 i1356_3_lut (.A(\mem[8] [6]), .B(\mem[9] [6]), .C(address[0]), 
         .Z(n1426)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1356_3_lut.init = 16'hcaca;
    LUT4 i1520_3_lut (.A(\mem[58] [0]), .B(\mem[59] [0]), .C(address[0]), 
         .Z(n1590)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1520_3_lut.init = 16'hcaca;
    LUT4 i1235_3_lut (.A(\mem[14] [1]), .B(\mem[15] [1]), .C(address[0]), 
         .Z(n1305)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1235_3_lut.init = 16'hcaca;
    LUT4 i1234_3_lut (.A(\mem[12] [1]), .B(\mem[13] [1]), .C(address[0]), 
         .Z(n1304)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1234_3_lut.init = 16'hcaca;
    LUT4 i1233_3_lut (.A(\mem[10] [1]), .B(\mem[11] [1]), .C(address[0]), 
         .Z(n1303)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1233_3_lut.init = 16'hcaca;
    LUT4 i1232_3_lut (.A(\mem[8] [1]), .B(\mem[9] [1]), .C(address[0]), 
         .Z(n1302)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1232_3_lut.init = 16'hcaca;
    LUT4 i1231_3_lut (.A(\mem[6] [1]), .B(\mem[7] [1]), .C(address[0]), 
         .Z(n1301)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1231_3_lut.init = 16'hcaca;
    LUT4 i1230_3_lut (.A(\mem[4] [1]), .B(\mem[5] [1]), .C(address[0]), 
         .Z(n1300)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1230_3_lut.init = 16'hcaca;
    PFUMX i1432 (.BLUT(n1488), .ALUT(n1489), .C0(address[1]), .Z(n1502));
    LUT4 i1243_3_lut (.A(\mem[30] [1]), .B(\mem[31] [1]), .C(address[0]), 
         .Z(n1313)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1243_3_lut.init = 16'hcaca;
    LUT4 i1242_3_lut (.A(\mem[28] [1]), .B(\mem[29] [1]), .C(address[0]), 
         .Z(n1312)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1242_3_lut.init = 16'hcaca;
    LUT4 i1663_3_lut (.A(\mem[34] [5]), .B(\mem[35] [5]), .C(address[0]), 
         .Z(n1733)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1663_3_lut.init = 16'hcaca;
    LUT4 i1229_3_lut (.A(\mem[2] [1]), .B(\mem[3] [1]), .C(address[0]), 
         .Z(n1299)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1229_3_lut.init = 16'hcaca;
    LUT4 i1228_3_lut (.A(\mem[0] [1]), .B(\mem[1] [1]), .C(address[0]), 
         .Z(n1298)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1228_3_lut.init = 16'hcaca;
    LUT4 i1700_3_lut (.A(\mem[46] [1]), .B(\mem[47] [1]), .C(address[0]), 
         .Z(n1770)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1700_3_lut.init = 16'hcaca;
    LUT4 i1646_3_lut (.A(\mem[62] [4]), .B(\mem[63] [4]), .C(address[0]), 
         .Z(n1716)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1646_3_lut.init = 16'hcaca;
    LUT4 i1521_3_lut (.A(\mem[60] [0]), .B(\mem[61] [0]), .C(address[0]), 
         .Z(n1591)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1521_3_lut.init = 16'hcaca;
    LUT4 i1662_3_lut (.A(\mem[32] [5]), .B(\mem[33] [5]), .C(address[0]), 
         .Z(n1732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1662_3_lut.init = 16'hcaca;
    LUT4 i1645_3_lut (.A(\mem[60] [4]), .B(\mem[61] [4]), .C(address[0]), 
         .Z(n1715)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1645_3_lut.init = 16'hcaca;
    LUT4 i1389_3_lut (.A(\mem[12] [2]), .B(\mem[13] [2]), .C(address[0]), 
         .Z(n1459)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1389_3_lut.init = 16'hcaca;
    LUT4 i1644_3_lut (.A(\mem[58] [4]), .B(\mem[59] [4]), .C(address[0]), 
         .Z(n1714)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1644_3_lut.init = 16'hcaca;
    LUT4 i1386_3_lut (.A(\mem[6] [2]), .B(\mem[7] [2]), .C(address[0]), 
         .Z(n1456)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1386_3_lut.init = 16'hcaca;
    LUT4 i1390_3_lut (.A(\mem[14] [2]), .B(\mem[15] [2]), .C(address[0]), 
         .Z(n1460)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1390_3_lut.init = 16'hcaca;
    LUT4 i1643_3_lut (.A(\mem[56] [4]), .B(\mem[57] [4]), .C(address[0]), 
         .Z(n1713)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1643_3_lut.init = 16'hcaca;
    LUT4 i1699_3_lut (.A(\mem[44] [1]), .B(\mem[45] [1]), .C(address[0]), 
         .Z(n1769)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1699_3_lut.init = 16'hcaca;
    LUT4 i1522_3_lut (.A(\mem[62] [0]), .B(\mem[63] [0]), .C(address[0]), 
         .Z(n1592)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1522_3_lut.init = 16'hcaca;
    LUT4 i1355_3_lut (.A(\mem[6] [6]), .B(\mem[7] [6]), .C(address[0]), 
         .Z(n1425)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1355_3_lut.init = 16'hcaca;
    LUT4 i1457_3_lut (.A(\mem[24] [7]), .B(\mem[25] [7]), .C(address[0]), 
         .Z(n1527)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1457_3_lut.init = 16'hcaca;
    LUT4 i1354_3_lut (.A(\mem[4] [6]), .B(\mem[5] [6]), .C(address[0]), 
         .Z(n1424)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1354_3_lut.init = 16'hcaca;
    LUT4 i1642_3_lut (.A(\mem[54] [4]), .B(\mem[55] [4]), .C(address[0]), 
         .Z(n1712)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1642_3_lut.init = 16'hcaca;
    LUT4 i1397_3_lut (.A(\mem[28] [2]), .B(\mem[29] [2]), .C(address[0]), 
         .Z(n1467)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1397_3_lut.init = 16'hcaca;
    LUT4 i1641_3_lut (.A(\mem[52] [4]), .B(\mem[53] [4]), .C(address[0]), 
         .Z(n1711)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1641_3_lut.init = 16'hcaca;
    LUT4 i1448_3_lut (.A(\mem[6] [7]), .B(\mem[7] [7]), .C(address[0]), 
         .Z(n1518)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1448_3_lut.init = 16'hcaca;
    LUT4 i1398_3_lut (.A(\mem[30] [2]), .B(\mem[31] [2]), .C(address[0]), 
         .Z(n1468)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1398_3_lut.init = 16'hcaca;
    LUT4 i1387_3_lut (.A(\mem[8] [2]), .B(\mem[9] [2]), .C(address[0]), 
         .Z(n1457)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1387_3_lut.init = 16'hcaca;
    LUT4 i1553_3_lut (.A(\mem[62] [2]), .B(\mem[63] [2]), .C(address[0]), 
         .Z(n1623)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1553_3_lut.init = 16'hcaca;
    LUT4 i1456_3_lut (.A(\mem[22] [7]), .B(\mem[23] [7]), .C(address[0]), 
         .Z(n1526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1456_3_lut.init = 16'hcaca;
    LUT4 i1552_3_lut (.A(\mem[60] [2]), .B(\mem[61] [2]), .C(address[0]), 
         .Z(n1622)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1552_3_lut.init = 16'hcaca;
    LUT4 i1551_3_lut (.A(\mem[58] [2]), .B(\mem[59] [2]), .C(address[0]), 
         .Z(n1621)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1551_3_lut.init = 16'hcaca;
    LUT4 i1388_3_lut (.A(\mem[10] [2]), .B(\mem[11] [2]), .C(address[0]), 
         .Z(n1458)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1388_3_lut.init = 16'hcaca;
    LUT4 i1550_3_lut (.A(\mem[56] [2]), .B(\mem[57] [2]), .C(address[0]), 
         .Z(n1620)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1550_3_lut.init = 16'hcaca;
    LUT4 i1395_3_lut (.A(\mem[24] [2]), .B(\mem[25] [2]), .C(address[0]), 
         .Z(n1465)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1395_3_lut.init = 16'hcaca;
    LUT4 i1455_3_lut (.A(\mem[20] [7]), .B(\mem[21] [7]), .C(address[0]), 
         .Z(n1525)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1455_3_lut.init = 16'hcaca;
    LUT4 i1353_3_lut (.A(\mem[2] [6]), .B(\mem[3] [6]), .C(address[0]), 
         .Z(n1423)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1353_3_lut.init = 16'hcaca;
    LUT4 i1396_3_lut (.A(\mem[26] [2]), .B(\mem[27] [2]), .C(address[0]), 
         .Z(n1466)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1396_3_lut.init = 16'hcaca;
    LUT4 i1515_3_lut (.A(\mem[48] [0]), .B(\mem[49] [0]), .C(address[0]), 
         .Z(n1585)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1515_3_lut.init = 16'hcaca;
    LUT4 i1352_3_lut (.A(\mem[0] [6]), .B(\mem[1] [6]), .C(address[0]), 
         .Z(n1422)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1352_3_lut.init = 16'hcaca;
    LUT4 i1454_3_lut (.A(\mem[18] [7]), .B(\mem[19] [7]), .C(address[0]), 
         .Z(n1524)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1454_3_lut.init = 16'hcaca;
    LUT4 i1453_3_lut (.A(\mem[16] [7]), .B(\mem[17] [7]), .C(address[0]), 
         .Z(n1523)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1453_3_lut.init = 16'hcaca;
    LUT4 i1393_3_lut (.A(\mem[20] [2]), .B(\mem[21] [2]), .C(address[0]), 
         .Z(n1463)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1393_3_lut.init = 16'hcaca;
    LUT4 i1394_3_lut (.A(\mem[22] [2]), .B(\mem[23] [2]), .C(address[0]), 
         .Z(n1464)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1394_3_lut.init = 16'hcaca;
    LUT4 i1516_3_lut (.A(\mem[50] [0]), .B(\mem[51] [0]), .C(address[0]), 
         .Z(n1586)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1516_3_lut.init = 16'hcaca;
    LUT4 i1385_3_lut (.A(\mem[4] [2]), .B(\mem[5] [2]), .C(address[0]), 
         .Z(n1455)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1385_3_lut.init = 16'hcaca;
    PFUMX i1433 (.BLUT(n1490), .ALUT(n1491), .C0(address[1]), .Z(n1503));
    LUT4 i1545_3_lut (.A(\mem[46] [2]), .B(\mem[47] [2]), .C(address[0]), 
         .Z(n1615)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1545_3_lut.init = 16'hcaca;
    LUT4 i1549_3_lut (.A(\mem[54] [2]), .B(\mem[55] [2]), .C(address[0]), 
         .Z(n1619)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1549_3_lut.init = 16'hcaca;
    LUT4 i1391_3_lut (.A(\mem[16] [2]), .B(\mem[17] [2]), .C(address[0]), 
         .Z(n1461)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1391_3_lut.init = 16'hcaca;
    LUT4 i1517_3_lut (.A(\mem[52] [0]), .B(\mem[53] [0]), .C(address[0]), 
         .Z(n1587)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1517_3_lut.init = 16'hcaca;
    LUT4 i1548_3_lut (.A(\mem[52] [2]), .B(\mem[53] [2]), .C(address[0]), 
         .Z(n1618)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1548_3_lut.init = 16'hcaca;
    PFUMX i1589 (.BLUT(n1647), .ALUT(n1648), .C0(address[1]), .Z(n1659));
    LUT4 i1639_3_lut (.A(\mem[48] [4]), .B(\mem[49] [4]), .C(address[0]), 
         .Z(n1709)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1639_3_lut.init = 16'hcaca;
    LUT4 i1640_3_lut (.A(\mem[50] [4]), .B(\mem[51] [4]), .C(address[0]), 
         .Z(n1710)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1640_3_lut.init = 16'hcaca;
    LUT4 i1546_3_lut (.A(\mem[48] [2]), .B(\mem[49] [2]), .C(address[0]), 
         .Z(n1616)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1546_3_lut.init = 16'hcaca;
    LUT4 i1544_3_lut (.A(\mem[44] [2]), .B(\mem[45] [2]), .C(address[0]), 
         .Z(n1614)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1544_3_lut.init = 16'hcaca;
    LUT4 i1543_3_lut (.A(\mem[42] [2]), .B(\mem[43] [2]), .C(address[0]), 
         .Z(n1613)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1543_3_lut.init = 16'hcaca;
    PFUMX i1434 (.BLUT(n1492), .ALUT(n1493), .C0(address[1]), .Z(n1504));
    LUT4 i1542_3_lut (.A(\mem[40] [2]), .B(\mem[41] [2]), .C(address[0]), 
         .Z(n1612)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1542_3_lut.init = 16'hcaca;
    LUT4 i1638_3_lut (.A(\mem[46] [4]), .B(\mem[47] [4]), .C(address[0]), 
         .Z(n1708)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1638_3_lut.init = 16'hcaca;
    LUT4 i1547_3_lut (.A(\mem[50] [2]), .B(\mem[51] [2]), .C(address[0]), 
         .Z(n1617)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1547_3_lut.init = 16'hcaca;
    LUT4 i1637_3_lut (.A(\mem[44] [4]), .B(\mem[45] [4]), .C(address[0]), 
         .Z(n1707)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1637_3_lut.init = 16'hcaca;
    LUT4 i1636_3_lut (.A(\mem[42] [4]), .B(\mem[43] [4]), .C(address[0]), 
         .Z(n1706)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1636_3_lut.init = 16'hcaca;
    LUT4 i1635_3_lut (.A(\mem[40] [4]), .B(\mem[41] [4]), .C(address[0]), 
         .Z(n1705)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1635_3_lut.init = 16'hcaca;
    LUT4 i1541_3_lut (.A(\mem[38] [2]), .B(\mem[39] [2]), .C(address[0]), 
         .Z(n1611)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1541_3_lut.init = 16'hcaca;
    LUT4 i1540_3_lut (.A(\mem[36] [2]), .B(\mem[37] [2]), .C(address[0]), 
         .Z(n1610)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1540_3_lut.init = 16'hcaca;
    LUT4 i1384_3_lut (.A(\mem[2] [2]), .B(\mem[3] [2]), .C(address[0]), 
         .Z(n1454)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1384_3_lut.init = 16'hcaca;
    LUT4 i1539_3_lut (.A(\mem[34] [2]), .B(\mem[35] [2]), .C(address[0]), 
         .Z(n1609)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1539_3_lut.init = 16'hcaca;
    LUT4 i1538_3_lut (.A(\mem[32] [2]), .B(\mem[33] [2]), .C(address[0]), 
         .Z(n1608)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1538_3_lut.init = 16'hcaca;
    LUT4 i1238_3_lut (.A(\mem[20] [1]), .B(\mem[21] [1]), .C(address[0]), 
         .Z(n1308)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1238_3_lut.init = 16'hcaca;
    LUT4 i1634_3_lut (.A(\mem[38] [4]), .B(\mem[39] [4]), .C(address[0]), 
         .Z(n1704)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1634_3_lut.init = 16'hcaca;
    LUT4 i1633_3_lut (.A(\mem[36] [4]), .B(\mem[37] [4]), .C(address[0]), 
         .Z(n1703)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1633_3_lut.init = 16'hcaca;
    LUT4 i1698_3_lut (.A(\mem[42] [1]), .B(\mem[43] [1]), .C(address[0]), 
         .Z(n1768)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1698_3_lut.init = 16'hcaca;
    PFUMX i1435 (.BLUT(n1494), .ALUT(n1495), .C0(address[1]), .Z(n1505));
    LUT4 i1632_3_lut (.A(\mem[34] [4]), .B(\mem[35] [4]), .C(address[0]), 
         .Z(n1702)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1632_3_lut.init = 16'hcaca;
    LUT4 i1631_3_lut (.A(\mem[32] [4]), .B(\mem[33] [4]), .C(address[0]), 
         .Z(n1701)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1631_3_lut.init = 16'hcaca;
    PFUMX i1590 (.BLUT(n1649), .ALUT(n1650), .C0(address[1]), .Z(n1660));
    PFUMX i1436 (.BLUT(n1496), .ALUT(n1497), .C0(address[1]), .Z(n1506));
    PFUMX i1437 (.BLUT(n1498), .ALUT(n1499), .C0(address[1]), .Z(n1507));
    PFUMX i1591 (.BLUT(n1651), .ALUT(n1652), .C0(address[1]), .Z(n1661));
    PFUMX i1710 (.BLUT(n1765), .ALUT(n1766), .C0(address[1]), .Z(n1780));
    PFUMX i1468 (.BLUT(n1529), .ALUT(n1530), .C0(address[1]), .Z(n1538));
    LUT4 i1239_3_lut (.A(\mem[22] [1]), .B(\mem[23] [1]), .C(address[0]), 
         .Z(n1309)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1239_3_lut.init = 16'hcaca;
    PFUMX i1463 (.BLUT(n1519), .ALUT(n1520), .C0(address[1]), .Z(n1533));
    PFUMX i1711 (.BLUT(n1767), .ALUT(n1768), .C0(address[1]), .Z(n1781));
    PFUMX i1464 (.BLUT(n1521), .ALUT(n1522), .C0(address[1]), .Z(n1534));
    PFUMX i1465 (.BLUT(n1523), .ALUT(n1524), .C0(address[1]), .Z(n1535));
    PFUMX i1592 (.BLUT(n1653), .ALUT(n1654), .C0(address[1]), .Z(n1662));
    PFUMX i1250 (.BLUT(n1310), .ALUT(n1311), .C0(address[1]), .Z(n1320));
    PFUMX i1709 (.BLUT(n1763), .ALUT(n1764), .C0(address[1]), .Z(n1779));
    PFUMX i1461 (.BLUT(n1515), .ALUT(n1516), .C0(address[1]), .Z(n1531));
    PFUMX i1462 (.BLUT(n1517), .ALUT(n1518), .C0(address[1]), .Z(n1532));
    PFUMX i1399 (.BLUT(n1453), .ALUT(n1454), .C0(address[1]), .Z(n1469));
    PFUMX i1527 (.BLUT(n1585), .ALUT(n1586), .C0(address[1]), .Z(n1597));
    PFUMX i1526 (.BLUT(n1583), .ALUT(n1584), .C0(address[1]), .Z(n1596));
    PFUMX i1344 (.BLUT(n1405), .ALUT(n1406), .C0(address[1]), .Z(n1414));
    PFUMX i1343 (.BLUT(n1403), .ALUT(n1404), .C0(address[1]), .Z(n1413));
    PFUMX i1342 (.BLUT(n1401), .ALUT(n1402), .C0(address[1]), .Z(n1412));
    PFUMX i1525 (.BLUT(n1581), .ALUT(n1582), .C0(address[1]), .Z(n1595));
    PFUMX i1524 (.BLUT(n1579), .ALUT(n1580), .C0(address[1]), .Z(n1594));
    PFUMX i1341 (.BLUT(n1399), .ALUT(n1400), .C0(address[1]), .Z(n1411));
    PFUMX i1340 (.BLUT(n1397), .ALUT(n1398), .C0(address[1]), .Z(n1410));
    PFUMX i1339 (.BLUT(n1395), .ALUT(n1396), .C0(address[1]), .Z(n1409));
    PFUMX i1523 (.BLUT(n1577), .ALUT(n1578), .C0(address[1]), .Z(n1593));
    PFUMX i1338 (.BLUT(n1393), .ALUT(n1394), .C0(address[1]), .Z(n1408));
    PFUMX i1337 (.BLUT(n1391), .ALUT(n1392), .C0(address[1]), .Z(n1407));
    PFUMX i1716 (.BLUT(n1777), .ALUT(n1778), .C0(address[1]), .Z(n1786));
    PFUMX i1715 (.BLUT(n1775), .ALUT(n1776), .C0(address[1]), .Z(n1785));
    PFUMX i1685 (.BLUT(n1746), .ALUT(n1747), .C0(address[1]), .Z(n1755));
    PFUMX i1248 (.BLUT(n1306), .ALUT(n1307), .C0(address[1]), .Z(n1318));
    PFUMX i1714 (.BLUT(n1773), .ALUT(n1774), .C0(address[1]), .Z(n1784));
    PFUMX i1684 (.BLUT(n1744), .ALUT(n1745), .C0(address[1]), .Z(n1754));
    PFUMX i1623 (.BLUT(n1684), .ALUT(n1685), .C0(address[1]), .Z(n1693));
    PFUMX i1313 (.BLUT(n1374), .ALUT(n1375), .C0(address[1]), .Z(n1383));
    PFUMX i1312 (.BLUT(n1372), .ALUT(n1373), .C0(address[1]), .Z(n1382));
    PFUMX i1311 (.BLUT(n1370), .ALUT(n1371), .C0(address[1]), .Z(n1381));
    PFUMX i1310 (.BLUT(n1368), .ALUT(n1369), .C0(address[1]), .Z(n1380));
    PFUMX i1683 (.BLUT(n1742), .ALUT(n1743), .C0(address[1]), .Z(n1753));
    PFUMX i1622 (.BLUT(n1682), .ALUT(n1683), .C0(address[1]), .Z(n1692));
    PFUMX i1499 (.BLUT(n1560), .ALUT(n1561), .C0(address[1]), .Z(n1569));
    PFUMX i1309 (.BLUT(n1366), .ALUT(n1367), .C0(address[1]), .Z(n1379));
    PFUMX i1308 (.BLUT(n1364), .ALUT(n1365), .C0(address[1]), .Z(n1378));
    PFUMX i1621 (.BLUT(n1680), .ALUT(n1681), .C0(address[1]), .Z(n1691));
    PFUMX i1498 (.BLUT(n1558), .ALUT(n1559), .C0(address[1]), .Z(n1568));
    PFUMX i1307 (.BLUT(n1362), .ALUT(n1363), .C0(address[1]), .Z(n1377));
    PFUMX i1497 (.BLUT(n1556), .ALUT(n1557), .C0(address[1]), .Z(n1567));
    PFUMX i1306 (.BLUT(n1360), .ALUT(n1361), .C0(address[1]), .Z(n1376));
    PFUMX i1682 (.BLUT(n1740), .ALUT(n1741), .C0(address[1]), .Z(n1752));
    PFUMX i1620 (.BLUT(n1678), .ALUT(n1679), .C0(address[1]), .Z(n1690));
    PFUMX i1496 (.BLUT(n1554), .ALUT(n1555), .C0(address[1]), .Z(n1566));
    PFUMX i1495 (.BLUT(n1552), .ALUT(n1553), .C0(address[1]), .Z(n1565));
    PFUMX i1619 (.BLUT(n1676), .ALUT(n1677), .C0(address[1]), .Z(n1689));
    PFUMX i1494 (.BLUT(n1550), .ALUT(n1551), .C0(address[1]), .Z(n1564));
    PFUMX i1493 (.BLUT(n1548), .ALUT(n1549), .C0(address[1]), .Z(n1563));
    PFUMX i1713 (.BLUT(n1771), .ALUT(n1772), .C0(address[1]), .Z(n1783));
    PFUMX i1681 (.BLUT(n1738), .ALUT(n1739), .C0(address[1]), .Z(n1751));
    PFUMX i1618 (.BLUT(n1674), .ALUT(n1675), .C0(address[1]), .Z(n1688));
    PFUMX i1492 (.BLUT(n1546), .ALUT(n1547), .C0(address[1]), .Z(n1562));
    PFUMX i1617 (.BLUT(n1672), .ALUT(n1673), .C0(address[1]), .Z(n1687));
    PFUMX i1616 (.BLUT(n1670), .ALUT(n1671), .C0(address[1]), .Z(n1686));
    PFUMX i1680 (.BLUT(n1736), .ALUT(n1737), .C0(address[1]), .Z(n1750));
    PFUMX i1282 (.BLUT(n1343), .ALUT(n1344), .C0(address[1]), .Z(n1352));
    PFUMX i1281 (.BLUT(n1341), .ALUT(n1342), .C0(address[1]), .Z(n1351));
    PFUMX i1280 (.BLUT(n1339), .ALUT(n1340), .C0(address[1]), .Z(n1350));
    PFUMX i1279 (.BLUT(n1337), .ALUT(n1338), .C0(address[1]), .Z(n1349));
    PFUMX i1278 (.BLUT(n1335), .ALUT(n1336), .C0(address[1]), .Z(n1348));
    PFUMX i1277 (.BLUT(n1333), .ALUT(n1334), .C0(address[1]), .Z(n1347));
    PFUMX i1276 (.BLUT(n1331), .ALUT(n1332), .C0(address[1]), .Z(n1346));
    PFUMX i1275 (.BLUT(n1329), .ALUT(n1330), .C0(address[1]), .Z(n1345));
    L6MUX21 i1472 (.D0(n1537), .D1(n1538), .SD(address[2]), .Z(n1542));
    L6MUX21 i1471 (.D0(n1535), .D1(n1536), .SD(address[2]), .Z(n1541));
    L6MUX21 i1470 (.D0(n1533), .D1(n1534), .SD(address[2]), .Z(n1540));
    L6MUX21 i1469 (.D0(n1531), .D1(n1532), .SD(address[2]), .Z(n1539));
    L6MUX21 i1596 (.D0(n1661), .D1(n1662), .SD(address[2]), .Z(n1666));
    L6MUX21 i1595 (.D0(n1659), .D1(n1660), .SD(address[2]), .Z(n1665));
    L6MUX21 i1594 (.D0(n1657), .D1(n1658), .SD(address[2]), .Z(n1664));
    L6MUX21 i1593 (.D0(n1655), .D1(n1656), .SD(address[2]), .Z(n1663));
    L6MUX21 i1441 (.D0(n1506), .D1(n1507), .SD(address[2]), .Z(n1511));
    L6MUX21 i1440 (.D0(n1504), .D1(n1505), .SD(address[2]), .Z(n1510));
    L6MUX21 i1439 (.D0(n1502), .D1(n1503), .SD(address[2]), .Z(n1509));
    L6MUX21 i1438 (.D0(n1500), .D1(n1501), .SD(address[2]), .Z(n1508));
    L6MUX21 i1379 (.D0(n1444), .D1(n1445), .SD(address[2]), .Z(n1449));
    L6MUX21 i1378 (.D0(n1442), .D1(n1443), .SD(address[2]), .Z(n1448));
    L6MUX21 i1377 (.D0(n1440), .D1(n1441), .SD(address[2]), .Z(n1447));
    L6MUX21 i1376 (.D0(n1438), .D1(n1439), .SD(address[2]), .Z(n1446));
    L6MUX21 i1255 (.D0(n1320), .D1(n1321), .SD(address[2]), .Z(n1325));
    L6MUX21 i1658 (.D0(n1723), .D1(n1724), .SD(address[2]), .Z(n1728));
    L6MUX21 i1657 (.D0(n1721), .D1(n1722), .SD(address[2]), .Z(n1727));
    L6MUX21 i1254 (.D0(n1318), .D1(n1319), .SD(address[2]), .Z(n1324));
    L6MUX21 i1253 (.D0(n1316), .D1(n1317), .SD(address[2]), .Z(n1323));
    L6MUX21 i1252 (.D0(n1314), .D1(n1315), .SD(address[2]), .Z(n1322));
    L6MUX21 i1656 (.D0(n1719), .D1(n1720), .SD(address[2]), .Z(n1726));
    L6MUX21 i1655 (.D0(n1717), .D1(n1718), .SD(address[2]), .Z(n1725));
    L6MUX21 i1565 (.D0(n1630), .D1(n1631), .SD(address[2]), .Z(n1635));
    L6MUX21 i1564 (.D0(n1628), .D1(n1629), .SD(address[2]), .Z(n1634));
    L6MUX21 i1563 (.D0(n1626), .D1(n1627), .SD(address[2]), .Z(n1633));
    L6MUX21 i1562 (.D0(n1624), .D1(n1625), .SD(address[2]), .Z(n1632));
    L6MUX21 i1720 (.D0(n1785), .D1(n1786), .SD(address[2]), .Z(n1790));
    L6MUX21 i1719 (.D0(n1783), .D1(n1784), .SD(address[2]), .Z(n1789));
    L6MUX21 i1407 (.D0(n1469), .D1(n1470), .SD(address[2]), .Z(n1477));
    L6MUX21 i1408 (.D0(n1471), .D1(n1472), .SD(address[2]), .Z(n1478));
    L6MUX21 i1409 (.D0(n1473), .D1(n1474), .SD(address[2]), .Z(n1479));
    L6MUX21 i1410 (.D0(n1475), .D1(n1476), .SD(address[2]), .Z(n1480));
    L6MUX21 i1534 (.D0(n1599), .D1(n1600), .SD(address[2]), .Z(n1604));
    L6MUX21 i1533 (.D0(n1597), .D1(n1598), .SD(address[2]), .Z(n1603));
    L6MUX21 i1532 (.D0(n1595), .D1(n1596), .SD(address[2]), .Z(n1602));
    L6MUX21 i1531 (.D0(n1593), .D1(n1594), .SD(address[2]), .Z(n1601));
    L6MUX21 i1718 (.D0(n1781), .D1(n1782), .SD(address[2]), .Z(n1788));
    L6MUX21 i1717 (.D0(n1779), .D1(n1780), .SD(address[2]), .Z(n1787));
    L6MUX21 i1348 (.D0(n1413), .D1(n1414), .SD(address[2]), .Z(n1418));
    L6MUX21 i1347 (.D0(n1411), .D1(n1412), .SD(address[2]), .Z(n1417));
    L6MUX21 i1346 (.D0(n1409), .D1(n1410), .SD(address[2]), .Z(n1416));
    L6MUX21 i1345 (.D0(n1407), .D1(n1408), .SD(address[2]), .Z(n1415));
    L6MUX21 i1689 (.D0(n1754), .D1(n1755), .SD(address[2]), .Z(n1759));
    L6MUX21 i1688 (.D0(n1752), .D1(n1753), .SD(address[2]), .Z(n1758));
    L6MUX21 i1687 (.D0(n1750), .D1(n1751), .SD(address[2]), .Z(n1757));
    L6MUX21 i1317 (.D0(n1382), .D1(n1383), .SD(address[2]), .Z(n1387));
    L6MUX21 i1316 (.D0(n1380), .D1(n1381), .SD(address[2]), .Z(n1386));
    L6MUX21 i1315 (.D0(n1378), .D1(n1379), .SD(address[2]), .Z(n1385));
    L6MUX21 i1686 (.D0(n1748), .D1(n1749), .SD(address[2]), .Z(n1756));
    L6MUX21 i1627 (.D0(n1692), .D1(n1693), .SD(address[2]), .Z(n1697));
    L6MUX21 i1626 (.D0(n1690), .D1(n1691), .SD(address[2]), .Z(n1696));
    L6MUX21 i1625 (.D0(n1688), .D1(n1689), .SD(address[2]), .Z(n1695));
    L6MUX21 i1624 (.D0(n1686), .D1(n1687), .SD(address[2]), .Z(n1694));
    L6MUX21 i1503 (.D0(n1568), .D1(n1569), .SD(address[2]), .Z(n1573));
    L6MUX21 i1502 (.D0(n1566), .D1(n1567), .SD(address[2]), .Z(n1572));
    L6MUX21 i1501 (.D0(n1564), .D1(n1565), .SD(address[2]), .Z(n1571));
    L6MUX21 i1314 (.D0(n1376), .D1(n1377), .SD(address[2]), .Z(n1384));
    L6MUX21 i1500 (.D0(n1562), .D1(n1563), .SD(address[2]), .Z(n1570));
    L6MUX21 i1286 (.D0(n1351), .D1(n1352), .SD(address[2]), .Z(n1356));
    L6MUX21 i1285 (.D0(n1349), .D1(n1350), .SD(address[2]), .Z(n1355));
    L6MUX21 i1284 (.D0(n1347), .D1(n1348), .SD(address[2]), .Z(n1354));
    L6MUX21 i1283 (.D0(n1345), .D1(n1346), .SD(address[2]), .Z(n1353));
    L6MUX21 i1474 (.D0(n1541), .D1(n1542), .SD(address[3]), .Z(n1544));
    L6MUX21 i1473 (.D0(n1539), .D1(n1540), .SD(address[3]), .Z(n1543));
    L6MUX21 i1598 (.D0(n1665), .D1(n1666), .SD(address[3]), .Z(n1668));
    L6MUX21 i1597 (.D0(n1663), .D1(n1664), .SD(address[3]), .Z(n1667));
    L6MUX21 i1443 (.D0(n1510), .D1(n1511), .SD(address[3]), .Z(n1513));
    L6MUX21 i1442 (.D0(n1508), .D1(n1509), .SD(address[3]), .Z(n1512));
    L6MUX21 i1381 (.D0(n1448), .D1(n1449), .SD(address[3]), .Z(n1451));
    L6MUX21 i1380 (.D0(n1446), .D1(n1447), .SD(address[3]), .Z(n1450));
    L6MUX21 i1660 (.D0(n1727), .D1(n1728), .SD(address[3]), .Z(n1730));
    L6MUX21 i1257 (.D0(n1324), .D1(n1325), .SD(address[3]), .Z(n1327));
    L6MUX21 i1256 (.D0(n1322), .D1(n1323), .SD(address[3]), .Z(n1326));
    L6MUX21 i1659 (.D0(n1725), .D1(n1726), .SD(address[3]), .Z(n1729));
    L6MUX21 i1567 (.D0(n1634), .D1(n1635), .SD(address[3]), .Z(n1637));
    L6MUX21 i1566 (.D0(n1632), .D1(n1633), .SD(address[3]), .Z(n1636));
    L6MUX21 i1722 (.D0(n1789), .D1(n1790), .SD(address[3]), .Z(n1792));
    L6MUX21 i1721 (.D0(n1787), .D1(n1788), .SD(address[3]), .Z(n1791));
    L6MUX21 i1411 (.D0(n1477), .D1(n1478), .SD(address[3]), .Z(n1481));
    L6MUX21 i1536 (.D0(n1603), .D1(n1604), .SD(address[3]), .Z(n1606));
    L6MUX21 i1412 (.D0(n1479), .D1(n1480), .SD(address[3]), .Z(n1482));
    L6MUX21 i1535 (.D0(n1601), .D1(n1602), .SD(address[3]), .Z(n1605));
    L6MUX21 i1691 (.D0(n1758), .D1(n1759), .SD(address[3]), .Z(n1761));
    L6MUX21 i1690 (.D0(n1756), .D1(n1757), .SD(address[3]), .Z(n1760));
    L6MUX21 i1350 (.D0(n1417), .D1(n1418), .SD(address[3]), .Z(n1420));
    L6MUX21 i1349 (.D0(n1415), .D1(n1416), .SD(address[3]), .Z(n1419));
    L6MUX21 i1629 (.D0(n1696), .D1(n1697), .SD(address[3]), .Z(n1699));
    L6MUX21 i1319 (.D0(n1386), .D1(n1387), .SD(address[3]), .Z(n1389));
    L6MUX21 i1318 (.D0(n1384), .D1(n1385), .SD(address[3]), .Z(n1388));
    L6MUX21 i1628 (.D0(n1694), .D1(n1695), .SD(address[3]), .Z(n1698));
    L6MUX21 i1505 (.D0(n1572), .D1(n1573), .SD(address[3]), .Z(n1575));
    L6MUX21 i1504 (.D0(n1570), .D1(n1571), .SD(address[3]), .Z(n1574));
    L6MUX21 i1288 (.D0(n1355), .D1(n1356), .SD(address[3]), .Z(n1358));
    L6MUX21 i1287 (.D0(n1353), .D1(n1354), .SD(address[3]), .Z(n1357));
    PFUMX i90911_i1 (.BLUT(n1328), .ALUT(n1793), .C0(address[5]), .Z(data_7__N_66[1]));
    PFUMX i91514_i1 (.BLUT(n1359), .ALUT(n1762), .C0(address[5]), .Z(data_7__N_66[5]));
    PFUMX i92117_i1 (.BLUT(n1390), .ALUT(n1731), .C0(address[5]), .Z(data_7__N_66[4]));
    PFUMX i92720_i1 (.BLUT(n1421), .ALUT(n1700), .C0(address[5]), .Z(data_7__N_66[3]));
    PFUMX i93323_i1 (.BLUT(n1452), .ALUT(n1669), .C0(address[5]), .Z(data_7__N_66[6]));
    PFUMX i93926_i1 (.BLUT(n1483), .ALUT(n1638), .C0(address[5]), .Z(data_7__N_66[2]));
    PFUMX i94529_i1 (.BLUT(n1514), .ALUT(n1607), .C0(address[5]), .Z(data_7__N_66[0]));
    PFUMX i95132_i1 (.BLUT(n1545), .ALUT(n1576), .C0(address[5]), .Z(data_7__N_66[7]));
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module CPU8BIT2
//

module CPU8BIT2 (akku_o_c_0, clk_c, reset_c, n1891, n1296, n1290, 
            mem_12__7__N_121, data_7__N_79, pc_5__N_30, n1287, n1289, 
            mem_6__7__N_103, n1286, n1272, mem_58__7__N_259, GND_net, 
            data, akku_o_c_6, akku_o_c_7, akku_o_c_4, akku_o_c_5, 
            akku_o_c_2, akku_o_c_3, akku_o_c_1, address, n1890, akku_o_c_8, 
            n1293, mem_59__7__N_262, mem_60__7__N_265, n681, mem_61__7__N_268, 
            mem_62__7__N_271, n1295, n1283, mem_48__7__N_229, n1292, 
            mem_49__7__N_232, mem_50__7__N_235, mem_51__7__N_238, mem_52__7__N_241, 
            mem_53__7__N_244, mem_54__7__N_247, n1260, mem_40__7__N_205, 
            mem_41__7__N_208, mem_42__7__N_211, mem_43__7__N_214, mem_44__7__N_217, 
            mem_45__7__N_220, mem_46__7__N_223, n1284, mem_32__7__N_181, 
            mem_33__7__N_184, mem_34__7__N_187, mem_35__7__N_190, mem_36__7__N_193, 
            mem_37__7__N_196, mem_38__7__N_199, n684, mem_24__7__N_157, 
            mem_25__7__N_160, mem_26__7__N_163, mem_27__7__N_166, mem_28__7__N_169, 
            mem_29__7__N_172, mem_30__7__N_175, n1261, mem_16__7__N_133, 
            mem_17__7__N_136, mem_18__7__N_139, mem_19__7__N_142, mem_20__7__N_145, 
            mem_21__7__N_148, mem_22__7__N_151, mem_8__7__N_109, mem_9__7__N_112, 
            mem_10__7__N_115, mem_5__7__N_100, mem_57__7__N_256, mem_56__7__N_253, 
            mem_4__7__N_97, mem_3__7__N_94, mem_2__7__N_91, mem_1__7__N_88, 
            mem_0__7__N_83, mem_14__7__N_127, mem_13__7__N_124, mem_11__7__N_118);
    output akku_o_c_0;
    input clk_c;
    input reset_c;
    output n1891;
    input n1296;
    input n1290;
    output mem_12__7__N_121;
    output data_7__N_79;
    input [5:0]pc_5__N_30;
    input n1287;
    input n1289;
    output mem_6__7__N_103;
    input n1286;
    input n1272;
    output mem_58__7__N_259;
    input GND_net;
    input [7:0]data;
    output akku_o_c_6;
    output akku_o_c_7;
    output akku_o_c_4;
    output akku_o_c_5;
    output akku_o_c_2;
    output akku_o_c_3;
    output akku_o_c_1;
    output [5:0]address;
    output n1890;
    output akku_o_c_8;
    input n1293;
    output mem_59__7__N_262;
    output mem_60__7__N_265;
    input n681;
    output mem_61__7__N_268;
    output mem_62__7__N_271;
    input n1295;
    input n1283;
    output mem_48__7__N_229;
    input n1292;
    output mem_49__7__N_232;
    output mem_50__7__N_235;
    output mem_51__7__N_238;
    output mem_52__7__N_241;
    output mem_53__7__N_244;
    output mem_54__7__N_247;
    input n1260;
    output mem_40__7__N_205;
    output mem_41__7__N_208;
    output mem_42__7__N_211;
    output mem_43__7__N_214;
    output mem_44__7__N_217;
    output mem_45__7__N_220;
    output mem_46__7__N_223;
    input n1284;
    output mem_32__7__N_181;
    output mem_33__7__N_184;
    output mem_34__7__N_187;
    output mem_35__7__N_190;
    output mem_36__7__N_193;
    output mem_37__7__N_196;
    output mem_38__7__N_199;
    input n684;
    output mem_24__7__N_157;
    output mem_25__7__N_160;
    output mem_26__7__N_163;
    output mem_27__7__N_166;
    output mem_28__7__N_169;
    output mem_29__7__N_172;
    output mem_30__7__N_175;
    input n1261;
    output mem_16__7__N_133;
    output mem_17__7__N_136;
    output mem_18__7__N_139;
    output mem_19__7__N_142;
    output mem_20__7__N_145;
    output mem_21__7__N_148;
    output mem_22__7__N_151;
    output mem_8__7__N_109;
    output mem_9__7__N_112;
    output mem_10__7__N_115;
    output mem_5__7__N_100;
    output mem_57__7__N_256;
    output mem_56__7__N_253;
    output mem_4__7__N_97;
    output mem_3__7__N_94;
    output mem_2__7__N_91;
    output mem_1__7__N_88;
    output mem_0__7__N_83;
    output mem_14__7__N_127;
    output mem_13__7__N_124;
    output mem_11__7__N_118;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(8[13:16])
    wire mem_12__7__N_121 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_12__7__N_121 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_6__7__N_103 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_6__7__N_103 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_58__7__N_259 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_58__7__N_259 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_59__7__N_262 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_59__7__N_262 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_60__7__N_265 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_60__7__N_265 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_61__7__N_268 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_61__7__N_268 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_62__7__N_271 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_62__7__N_271 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_48__7__N_229 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_48__7__N_229 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_49__7__N_232 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_49__7__N_232 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_50__7__N_235 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_50__7__N_235 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_51__7__N_238 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_51__7__N_238 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_52__7__N_241 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_52__7__N_241 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_53__7__N_244 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_53__7__N_244 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_54__7__N_247 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_54__7__N_247 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_40__7__N_205 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_40__7__N_205 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_41__7__N_208 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_41__7__N_208 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_42__7__N_211 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_42__7__N_211 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_43__7__N_214 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_43__7__N_214 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_44__7__N_217 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_44__7__N_217 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_45__7__N_220 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_45__7__N_220 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_46__7__N_223 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_46__7__N_223 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_32__7__N_181 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_32__7__N_181 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_33__7__N_184 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_33__7__N_184 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_34__7__N_187 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_34__7__N_187 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_35__7__N_190 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_35__7__N_190 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_36__7__N_193 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_36__7__N_193 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_37__7__N_196 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_37__7__N_196 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_38__7__N_199 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_38__7__N_199 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_24__7__N_157 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_24__7__N_157 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_25__7__N_160 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_25__7__N_160 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_26__7__N_163 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_26__7__N_163 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_27__7__N_166 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_27__7__N_166 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_28__7__N_169 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_28__7__N_169 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_29__7__N_172 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_29__7__N_172 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_30__7__N_175 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_30__7__N_175 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_16__7__N_133 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_16__7__N_133 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_17__7__N_136 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_17__7__N_136 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_18__7__N_139 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_18__7__N_139 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_19__7__N_142 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_19__7__N_142 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_20__7__N_145 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_20__7__N_145 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_21__7__N_148 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_21__7__N_148 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_22__7__N_151 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_22__7__N_151 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_8__7__N_109 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_8__7__N_109 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_9__7__N_112 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_9__7__N_112 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_10__7__N_115 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_10__7__N_115 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_5__7__N_100 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_5__7__N_100 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_57__7__N_256 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_57__7__N_256 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_56__7__N_253 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_56__7__N_253 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_4__7__N_97 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_4__7__N_97 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_3__7__N_94 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_3__7__N_94 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_2__7__N_91 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_2__7__N_91 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_1__7__N_88 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_1__7__N_88 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_0__7__N_83 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_0__7__N_83 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_14__7__N_127 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_14__7__N_127 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_13__7__N_124 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_13__7__N_124 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_11__7__N_118 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_11__7__N_118 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [2:0]states;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(25[15:21])
    
    wire clk_c_enable_7, clk_c_enable_15;
    wire [8:0]akku_o_8__N_44;
    
    wire n1979, n1895, n1889, n430, n2;
    wire [5:0]pc;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(23[15:17])
    wire [2:0]states_2__N_53;
    wire [5:0]pc_5__N_30_c;
    
    wire n1243, n1242;
    wire [7:0]akku_o_8__N_36;
    
    wire n1241, n1240, n1239, n1894, n1892, clk_c_enable_8;
    wire [8:0]akku_o_8__N_11;
    wire [5:0]adress_5__N_3;
    
    LUT4 i661_1_lut_3_lut (.A(states[1]), .B(states[2]), .C(states[0]), 
         .Z(clk_c_enable_7)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[33:48])
    defparam i661_1_lut_3_lut.init = 16'h0101;
    FD1P3AX akku_i1 (.D(akku_o_8__N_44[0]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_0)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam akku_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_81 (.A(reset_c), .B(clk_c), .Z(n1979)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_rep_81.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n1891), .B(n1979), .C(n1296), .D(n1290), 
         .Z(mem_12__7__N_121)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i1_3_lut_3_lut_2_lut_3_lut_4_lut (.A(reset_c), .B(clk_c), .C(states[0]), 
         .D(states[1]), .Z(data_7__N_79)) /* synthesis lut_function=(!((B+!((D)+!C))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_3_lut_3_lut_2_lut_3_lut_4_lut.init = 16'h2202;
    FD1S3IX states__i2 (.D(n1889), .CK(clk_c), .CD(n1895), .Q(states[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam states__i2.GSR = "ENABLED";
    FD1S3IX states__i1 (.D(n2), .CK(clk_c), .CD(n430), .Q(states[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam states__i1.GSR = "ENABLED";
    FD1P3AX pc_i0_i0 (.D(pc_5__N_30[0]), .SP(clk_c_enable_7), .CK(clk_c), 
            .Q(pc[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam pc_i0_i0.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_8 (.A(n1891), .B(n1979), .C(n1287), 
         .D(n1289), .Z(mem_6__7__N_103)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_8.init = 16'h0004;
    FD1S3IX states__i0 (.D(states_2__N_53[0]), .CK(clk_c), .CD(n1895), 
            .Q(states[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam states__i0.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_9 (.A(n1891), .B(n1979), .C(n1286), 
         .D(n1272), .Z(mem_58__7__N_259)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_9.init = 16'h0400;
    FD1P3AX pc_i0_i5 (.D(pc_5__N_30_c[5]), .SP(clk_c_enable_7), .CK(clk_c), 
            .Q(pc[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam pc_i0_i5.GSR = "ENABLED";
    CCU2D add_91_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n1243), 
          .S0(akku_o_8__N_44[8]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(47[39:69])
    defparam add_91_cout.INIT0 = 16'h0000;
    defparam add_91_cout.INIT1 = 16'h0000;
    defparam add_91_cout.INJECT1_0 = "NO";
    defparam add_91_cout.INJECT1_1 = "NO";
    CCU2D add_91_9 (.A0(data[6]), .B0(states[0]), .C0(akku_o_8__N_36[6]), 
          .D0(akku_o_c_6), .A1(data[7]), .B1(states[0]), .C1(akku_o_8__N_36[7]), 
          .D1(akku_o_c_7), .CIN(n1242), .COUT(n1243), .S0(akku_o_8__N_44[6]), 
          .S1(akku_o_8__N_44[7]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(47[39:69])
    defparam add_91_9.INIT0 = 16'hd1e2;
    defparam add_91_9.INIT1 = 16'hd1e2;
    defparam add_91_9.INJECT1_0 = "NO";
    defparam add_91_9.INJECT1_1 = "NO";
    CCU2D add_91_7 (.A0(data[4]), .B0(states[0]), .C0(akku_o_8__N_36[4]), 
          .D0(akku_o_c_4), .A1(data[5]), .B1(states[0]), .C1(akku_o_8__N_36[5]), 
          .D1(akku_o_c_5), .CIN(n1241), .COUT(n1242), .S0(akku_o_8__N_44[4]), 
          .S1(akku_o_8__N_44[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(47[39:69])
    defparam add_91_7.INIT0 = 16'hd1e2;
    defparam add_91_7.INIT1 = 16'hd1e2;
    defparam add_91_7.INJECT1_0 = "NO";
    defparam add_91_7.INJECT1_1 = "NO";
    CCU2D add_91_5 (.A0(data[2]), .B0(states[0]), .C0(akku_o_8__N_36[2]), 
          .D0(akku_o_c_2), .A1(data[3]), .B1(states[0]), .C1(akku_o_8__N_36[3]), 
          .D1(akku_o_c_3), .CIN(n1240), .COUT(n1241), .S0(akku_o_8__N_44[2]), 
          .S1(akku_o_8__N_44[3]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(47[39:69])
    defparam add_91_5.INIT0 = 16'hd1e2;
    defparam add_91_5.INIT1 = 16'hd1e2;
    defparam add_91_5.INJECT1_0 = "NO";
    defparam add_91_5.INJECT1_1 = "NO";
    CCU2D add_91_3 (.A0(data[0]), .B0(states[0]), .C0(akku_o_8__N_36[0]), 
          .D0(akku_o_c_0), .A1(data[1]), .B1(states[0]), .C1(akku_o_8__N_36[1]), 
          .D1(akku_o_c_1), .CIN(n1239), .COUT(n1240), .S0(akku_o_8__N_44[0]), 
          .S1(akku_o_8__N_44[1]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(47[39:69])
    defparam add_91_3.INIT0 = 16'hd1e2;
    defparam add_91_3.INIT1 = 16'hd1e2;
    defparam add_91_3.INJECT1_0 = "NO";
    defparam add_91_3.INJECT1_1 = "NO";
    LUT4 i132_2_lut_3_lut_4_lut (.A(address[2]), .B(n1894), .C(address[4]), 
         .D(address[3]), .Z(pc_5__N_30_c[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i132_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i1_2_lut_rep_73_3_lut_4_lut (.A(states[1]), .B(states[0]), .C(n1979), 
         .D(states[2]), .Z(n1890)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_rep_73_3_lut_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_rep_74_3_lut (.A(states[1]), .B(states[0]), .C(states[2]), 
         .Z(n1891)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_rep_74_3_lut.init = 16'hfbfb;
    LUT4 i113_2_lut_rep_77 (.A(address[1]), .B(address[0]), .Z(n1894)) /* synthesis lut_function=(A (B)) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i113_2_lut_rep_77.init = 16'h8888;
    LUT4 i120_2_lut_rep_75_3_lut (.A(address[1]), .B(address[0]), .C(address[2]), 
         .Z(n1892)) /* synthesis lut_function=(A (B (C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i120_2_lut_rep_75_3_lut.init = 16'h8080;
    LUT4 i385_2_lut_3_lut_4_lut (.A(data[7]), .B(akku_o_c_8), .C(n1895), 
         .D(data[6]), .Z(n430)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i385_2_lut_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_10 (.A(n1891), .B(n1979), .C(n1293), 
         .D(n1272), .Z(mem_59__7__N_262)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_10.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_11 (.A(n1891), .B(n1979), .C(n1296), 
         .D(n1272), .Z(mem_60__7__N_265)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_11.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_12 (.A(n1891), .B(n1979), .C(n681), 
         .D(n1272), .Z(mem_61__7__N_268)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_12.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_13 (.A(n1891), .B(n1979), .C(n1287), 
         .D(n1272), .Z(mem_62__7__N_271)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_13.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_14 (.A(n1891), .B(n1979), .C(n1295), 
         .D(n1283), .Z(mem_48__7__N_229)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_14.init = 16'h0004;
    LUT4 i366_2_lut_rep_80 (.A(states[1]), .B(states[2]), .Z(clk_c_enable_15)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(46[13] 52[22])
    defparam i366_2_lut_rep_80.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_4_lut_adj_15 (.A(n1891), .B(n1979), .C(n1292), 
         .D(n1283), .Z(mem_49__7__N_232)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_15.init = 16'h0004;
    LUT4 i13_4_lut_3_lut (.A(states[1]), .B(states[2]), .C(states[0]), 
         .Z(clk_c_enable_8)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(46[13] 52[22])
    defparam i13_4_lut_3_lut.init = 16'h4242;
    LUT4 i1_2_lut_3_lut_4_lut_adj_16 (.A(n1891), .B(n1979), .C(n1286), 
         .D(n1283), .Z(mem_50__7__N_235)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_16.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_17 (.A(n1891), .B(n1979), .C(n1293), 
         .D(n1283), .Z(mem_51__7__N_238)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_17.init = 16'h0004;
    LUT4 i118_2_lut_3_lut (.A(address[1]), .B(address[0]), .C(address[2]), 
         .Z(pc_5__N_30_c[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i118_2_lut_3_lut.init = 16'h7878;
    LUT4 i1_2_lut_3_lut_4_lut_adj_18 (.A(n1891), .B(n1979), .C(n1296), 
         .D(n1283), .Z(mem_52__7__N_241)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_18.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_19 (.A(n1891), .B(n1979), .C(n681), 
         .D(n1283), .Z(mem_53__7__N_244)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_19.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_20 (.A(n1891), .B(n1979), .C(n1287), 
         .D(n1283), .Z(mem_54__7__N_247)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_20.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_21 (.A(n1891), .B(n1979), .C(n1295), 
         .D(n1260), .Z(mem_40__7__N_205)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_21.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_22 (.A(n1891), .B(n1979), .C(n1292), 
         .D(n1260), .Z(mem_41__7__N_208)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_22.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_23 (.A(n1891), .B(n1979), .C(n1286), 
         .D(n1260), .Z(mem_42__7__N_211)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_23.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_24 (.A(n1891), .B(n1979), .C(n1293), 
         .D(n1260), .Z(mem_43__7__N_214)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_24.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_25 (.A(n1891), .B(n1979), .C(n1296), 
         .D(n1260), .Z(mem_44__7__N_217)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_25.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_26 (.A(n1891), .B(n1979), .C(n681), 
         .D(n1260), .Z(mem_45__7__N_220)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_26.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_27 (.A(n1891), .B(n1979), .C(n1287), 
         .D(n1260), .Z(mem_46__7__N_223)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_27.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_28 (.A(n1891), .B(n1979), .C(n1295), 
         .D(n1284), .Z(mem_32__7__N_181)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_28.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_29 (.A(n1891), .B(n1979), .C(n1292), 
         .D(n1284), .Z(mem_33__7__N_184)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_29.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_30 (.A(n1891), .B(n1979), .C(n1286), 
         .D(n1284), .Z(mem_34__7__N_187)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_30.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_31 (.A(n1891), .B(n1979), .C(n1293), 
         .D(n1284), .Z(mem_35__7__N_190)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_31.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_32 (.A(n1891), .B(n1979), .C(n1296), 
         .D(n1284), .Z(mem_36__7__N_193)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_32.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_33 (.A(n1891), .B(n1979), .C(n681), 
         .D(n1284), .Z(mem_37__7__N_196)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_33.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_34 (.A(n1891), .B(n1979), .C(n1287), 
         .D(n1284), .Z(mem_38__7__N_199)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_34.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_35 (.A(n1891), .B(n1979), .C(n1295), 
         .D(n684), .Z(mem_24__7__N_157)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_35.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_36 (.A(n1891), .B(n1979), .C(n1292), 
         .D(n684), .Z(mem_25__7__N_160)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_36.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_37 (.A(n1891), .B(n1979), .C(n1286), 
         .D(n684), .Z(mem_26__7__N_163)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_37.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_38 (.A(n1891), .B(n1979), .C(n1293), 
         .D(n684), .Z(mem_27__7__N_166)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_38.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_39 (.A(n1891), .B(n1979), .C(n1296), 
         .D(n684), .Z(mem_28__7__N_169)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_39.init = 16'h0004;
    LUT4 i125_2_lut_3_lut_4_lut (.A(address[1]), .B(address[0]), .C(address[3]), 
         .D(address[2]), .Z(pc_5__N_30_c[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i125_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_40 (.A(n1891), .B(n1979), .C(n681), 
         .D(n684), .Z(mem_29__7__N_172)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_40.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_41 (.A(n1891), .B(n1979), .C(n1287), 
         .D(n684), .Z(mem_30__7__N_175)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_41.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_42 (.A(n1891), .B(n1979), .C(n1295), 
         .D(n1261), .Z(mem_16__7__N_133)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_42.init = 16'h0004;
    LUT4 i1_2_lut_rep_72_3_lut (.A(data[7]), .B(akku_o_c_8), .C(data[6]), 
         .Z(n1889)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_72_3_lut.init = 16'h8080;
    LUT4 i885_2_lut_3_lut (.A(data[7]), .B(akku_o_c_8), .C(data[6]), .Z(states_2__N_53[0])) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;
    defparam i885_2_lut_3_lut.init = 16'h8f8f;
    LUT4 i2_3_lut_rep_78 (.A(states[1]), .B(states[2]), .C(states[0]), 
         .Z(n1895)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[33:48])
    defparam i2_3_lut_rep_78.init = 16'hfefe;
    LUT4 i145_1_lut (.A(data[7]), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(57[20:43])
    defparam i145_1_lut.init = 16'h5555;
    LUT4 i139_3_lut_4_lut (.A(address[3]), .B(n1892), .C(address[4]), 
         .D(address[5]), .Z(pc_5__N_30_c[5])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i139_3_lut_4_lut.init = 16'h7f80;
    FD1P3AX pc_i0_i4 (.D(pc_5__N_30_c[4]), .SP(clk_c_enable_7), .CK(clk_c), 
            .Q(pc[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam pc_i0_i4.GSR = "ENABLED";
    FD1P3AX pc_i0_i3 (.D(pc_5__N_30_c[3]), .SP(clk_c_enable_7), .CK(clk_c), 
            .Q(pc[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam pc_i0_i3.GSR = "ENABLED";
    FD1P3AX pc_i0_i2 (.D(pc_5__N_30_c[2]), .SP(clk_c_enable_7), .CK(clk_c), 
            .Q(pc[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam pc_i0_i2.GSR = "ENABLED";
    LUT4 i1968_2_lut (.A(akku_o_c_6), .B(data[6]), .Z(akku_o_8__N_36[6])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(49[60:94])
    defparam i1968_2_lut.init = 16'h1111;
    FD1P3AX pc_i0_i1 (.D(pc_5__N_30_c[1]), .SP(clk_c_enable_7), .CK(clk_c), 
            .Q(pc[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam pc_i0_i1.GSR = "ENABLED";
    FD1P3AX akku_i9 (.D(akku_o_8__N_11[8]), .SP(clk_c_enable_8), .CK(clk_c), 
            .Q(akku_o_c_8)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam akku_i9.GSR = "ENABLED";
    CCU2D add_91_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(states[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n1239));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(47[39:69])
    defparam add_91_1.INIT0 = 16'hF000;
    defparam add_91_1.INIT1 = 16'h0fff;
    defparam add_91_1.INJECT1_0 = "NO";
    defparam add_91_1.INJECT1_1 = "NO";
    LUT4 i1965_2_lut (.A(akku_o_c_7), .B(data[7]), .Z(akku_o_8__N_36[7])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(49[60:94])
    defparam i1965_2_lut.init = 16'h1111;
    LUT4 i1974_2_lut (.A(akku_o_c_4), .B(data[4]), .Z(akku_o_8__N_36[4])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(49[60:94])
    defparam i1974_2_lut.init = 16'h1111;
    LUT4 i1971_2_lut (.A(akku_o_c_5), .B(data[5]), .Z(akku_o_8__N_36[5])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(49[60:94])
    defparam i1971_2_lut.init = 16'h1111;
    FD1P3AX akku_i8 (.D(akku_o_8__N_44[7]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_7)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam akku_i8.GSR = "ENABLED";
    LUT4 i1980_2_lut (.A(akku_o_c_2), .B(data[2]), .Z(akku_o_8__N_36[2])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(49[60:94])
    defparam i1980_2_lut.init = 16'h1111;
    FD1P3AX akku_i7 (.D(akku_o_8__N_44[6]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_6)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam akku_i7.GSR = "ENABLED";
    FD1P3AX akku_i6 (.D(akku_o_8__N_44[5]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_5)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam akku_i6.GSR = "ENABLED";
    FD1P3AX akku_i5 (.D(akku_o_8__N_44[4]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_4)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam akku_i5.GSR = "ENABLED";
    FD1P3AX akku_i4 (.D(akku_o_8__N_44[3]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_3)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam akku_i4.GSR = "ENABLED";
    LUT4 i1977_2_lut (.A(akku_o_c_3), .B(data[3]), .Z(akku_o_8__N_36[3])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(49[60:94])
    defparam i1977_2_lut.init = 16'h1111;
    LUT4 i1962_2_lut (.A(akku_o_c_0), .B(data[0]), .Z(akku_o_8__N_36[0])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(49[60:94])
    defparam i1962_2_lut.init = 16'h1111;
    FD1P3AX akku_i3 (.D(akku_o_8__N_44[2]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_2)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam akku_i3.GSR = "ENABLED";
    FD1P3AX akku_i2 (.D(akku_o_8__N_44[1]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_1)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam akku_i2.GSR = "ENABLED";
    LUT4 i1959_2_lut (.A(akku_o_c_1), .B(data[1]), .Z(akku_o_8__N_36[1])) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(49[60:94])
    defparam i1959_2_lut.init = 16'h1111;
    FD1S3AX adreg_i5 (.D(adress_5__N_3[5]), .CK(clk_c), .Q(address[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam adreg_i5.GSR = "ENABLED";
    FD1S3AX adreg_i4 (.D(adress_5__N_3[4]), .CK(clk_c), .Q(address[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam adreg_i4.GSR = "ENABLED";
    FD1S3AX adreg_i3 (.D(adress_5__N_3[3]), .CK(clk_c), .Q(address[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam adreg_i3.GSR = "ENABLED";
    LUT4 i111_2_lut (.A(address[1]), .B(address[0]), .Z(pc_5__N_30_c[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i111_2_lut.init = 16'h6666;
    LUT4 i891_2_lut (.A(akku_o_8__N_44[8]), .B(states[2]), .Z(akku_o_8__N_11[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(46[13] 52[22])
    defparam i891_2_lut.init = 16'h2222;
    FD1S3AX adreg_i2 (.D(adress_5__N_3[2]), .CK(clk_c), .Q(address[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam adreg_i2.GSR = "ENABLED";
    FD1S3AX adreg_i1 (.D(adress_5__N_3[1]), .CK(clk_c), .Q(address[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam adreg_i1.GSR = "ENABLED";
    LUT4 pc_5__I_0_85_i6_3_lut (.A(data[5]), .B(pc[5]), .C(n1895), .Z(adress_5__N_3[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(36[13] 43[20])
    defparam pc_5__I_0_85_i6_3_lut.init = 16'hcaca;
    LUT4 pc_5__I_0_85_i5_3_lut (.A(data[4]), .B(pc[4]), .C(n1895), .Z(adress_5__N_3[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(36[13] 43[20])
    defparam pc_5__I_0_85_i5_3_lut.init = 16'hcaca;
    LUT4 pc_5__I_0_85_i4_3_lut (.A(data[3]), .B(pc[3]), .C(n1895), .Z(adress_5__N_3[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(36[13] 43[20])
    defparam pc_5__I_0_85_i4_3_lut.init = 16'hcaca;
    LUT4 pc_5__I_0_85_i3_3_lut (.A(data[2]), .B(pc[2]), .C(n1895), .Z(adress_5__N_3[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(36[13] 43[20])
    defparam pc_5__I_0_85_i3_3_lut.init = 16'hcaca;
    LUT4 pc_5__I_0_85_i2_3_lut (.A(data[1]), .B(pc[1]), .C(n1895), .Z(adress_5__N_3[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(36[13] 43[20])
    defparam pc_5__I_0_85_i2_3_lut.init = 16'hcaca;
    LUT4 pc_5__I_0_85_i1_3_lut (.A(data[0]), .B(pc[0]), .C(n1895), .Z(adress_5__N_3[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(36[13] 43[20])
    defparam pc_5__I_0_85_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_43 (.A(n1891), .B(n1979), .C(n1292), 
         .D(n1261), .Z(mem_17__7__N_136)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_43.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_44 (.A(n1891), .B(n1979), .C(n1286), 
         .D(n1261), .Z(mem_18__7__N_139)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_44.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_45 (.A(n1891), .B(n1979), .C(n1293), 
         .D(n1261), .Z(mem_19__7__N_142)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_45.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_46 (.A(n1891), .B(n1979), .C(n1296), 
         .D(n1261), .Z(mem_20__7__N_145)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_46.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_47 (.A(n1891), .B(n1979), .C(n681), 
         .D(n1261), .Z(mem_21__7__N_148)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_47.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_48 (.A(n1891), .B(n1979), .C(n1287), 
         .D(n1261), .Z(mem_22__7__N_151)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_48.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_49 (.A(n1891), .B(n1979), .C(n1295), 
         .D(n1290), .Z(mem_8__7__N_109)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_49.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_50 (.A(n1891), .B(n1979), .C(n1292), 
         .D(n1290), .Z(mem_9__7__N_112)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_50.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_51 (.A(n1891), .B(n1979), .C(n1286), 
         .D(n1290), .Z(mem_10__7__N_115)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_51.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_52 (.A(n1891), .B(n1979), .C(n681), 
         .D(n1289), .Z(mem_5__7__N_100)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_52.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_53 (.A(n1891), .B(n1979), .C(n1292), 
         .D(n1272), .Z(mem_57__7__N_256)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_53.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_54 (.A(n1891), .B(n1979), .C(n1295), 
         .D(n1272), .Z(mem_56__7__N_253)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_54.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_55 (.A(n1891), .B(n1979), .C(n1296), 
         .D(n1289), .Z(mem_4__7__N_97)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_55.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_56 (.A(n1891), .B(n1979), .C(n1293), 
         .D(n1289), .Z(mem_3__7__N_94)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_56.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_57 (.A(n1891), .B(n1979), .C(n1286), 
         .D(n1289), .Z(mem_2__7__N_91)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_57.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_58 (.A(n1891), .B(n1979), .C(n1292), 
         .D(n1289), .Z(mem_1__7__N_88)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_58.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_59 (.A(n1891), .B(n1979), .C(n1295), 
         .D(n1289), .Z(mem_0__7__N_83)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_59.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_60 (.A(n1891), .B(n1979), .C(n1287), 
         .D(n1290), .Z(mem_14__7__N_127)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_60.init = 16'h0004;
    FD1S3AX adreg_i0 (.D(adress_5__N_3[0]), .CK(clk_c), .Q(address[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 69[16])
    defparam adreg_i0.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_61 (.A(n1891), .B(n1979), .C(n681), 
         .D(n1290), .Z(mem_13__7__N_124)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_61.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_62 (.A(n1891), .B(n1979), .C(n1293), 
         .D(n1290), .Z(mem_11__7__N_118)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(80[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_62.init = 16'h0004;
    
endmodule
