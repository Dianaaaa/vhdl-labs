// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.11.0.396.4
// Netlist written on Fri Nov 20 10:28:22 2020
//
// Verilog Description of module cpu2system
//

module cpu2system (clk, reset, akku_o);   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(7[8:18])
    input clk;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(8[13:16])
    input reset;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(9[13:18])
    output [8:0]akku_o;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(8[13:16])
    wire mem_0__7__N_101 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_0__7__N_101 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_2__7__N_109 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_2__7__N_109 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_3__7__N_112 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_3__7__N_112 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_4__7__N_115 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_4__7__N_115 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_7__7__N_124 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_7__7__N_124 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_8__7__N_127 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_8__7__N_127 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_10__7__N_133 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_10__7__N_133 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_11__7__N_136 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_11__7__N_136 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_12__7__N_139 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_12__7__N_139 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_15__7__N_148 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_15__7__N_148 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_16__7__N_151 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_16__7__N_151 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_18__7__N_157 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_18__7__N_157 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_19__7__N_160 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_19__7__N_160 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_20__7__N_163 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_20__7__N_163 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_23__7__N_172 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_23__7__N_172 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_24__7__N_175 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_24__7__N_175 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_26__7__N_181 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_26__7__N_181 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_27__7__N_184 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_27__7__N_184 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_28__7__N_187 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_28__7__N_187 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_31__7__N_196 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_31__7__N_196 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_32__7__N_199 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_32__7__N_199 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_34__7__N_205 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_34__7__N_205 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_35__7__N_208 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_35__7__N_208 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_36__7__N_211 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_36__7__N_211 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_39__7__N_220 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_39__7__N_220 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_40__7__N_223 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_40__7__N_223 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_42__7__N_229 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_42__7__N_229 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_43__7__N_232 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_43__7__N_232 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_44__7__N_235 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_44__7__N_235 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_47__7__N_244 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_47__7__N_244 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_48__7__N_247 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_48__7__N_247 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_50__7__N_253 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_50__7__N_253 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_51__7__N_256 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_51__7__N_256 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_52__7__N_259 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_52__7__N_259 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_55__7__N_268 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_55__7__N_268 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_56__7__N_271 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_56__7__N_271 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_58__7__N_277 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_58__7__N_277 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_59__7__N_280 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_59__7__N_280 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_60__7__N_283 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_60__7__N_283 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_63__7__N_292 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_63__7__N_292 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire GND_net, reset_c, akku_o_c_8, akku_o_c_7, akku_o_c_6, akku_o_c_5, 
        akku_o_c_4, akku_o_c_3, akku_o_c_2, akku_o_c_1, akku_o_c_0;
    wire [7:0]data;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(37[13:17])
    wire [2:0]states_2__N_71;
    
    wire n1916, n1302;
    wire [5:0]address;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(24[9:16])
    
    wire n1911, data_7__N_97, n1910, n1327, n1906, n1905, n1902, 
        n1901, n1900, n1899, n1898, n1896, VCC_net, n1895, n1328;
    
    IB reset_pad (.I(reset), .O(reset_c));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(9[13:18])
    IB clk_pad (.I(clk), .O(clk_c));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(8[13:16])
    OB akku_o_pad_0 (.I(akku_o_c_0), .O(akku_o[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_1 (.I(akku_o_c_1), .O(akku_o[1]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_2 (.I(akku_o_c_2), .O(akku_o[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_3 (.I(akku_o_c_3), .O(akku_o[3]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_4 (.I(akku_o_c_4), .O(akku_o[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_5 (.I(akku_o_c_5), .O(akku_o[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_6 (.I(akku_o_c_6), .O(akku_o[6]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_7 (.I(akku_o_c_7), .O(akku_o[7]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_8 (.I(akku_o_c_8), .O(akku_o[8]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    VHI i1937 (.Z(VCC_net));
    VLO i1 (.Z(GND_net));
    TSALL TSALL_INST (.TSALL(GND_net));
    GSR GSR_INST (.GSR(reset_c));
    \sram64kx8("sram64kx8.dat")(1,13)  RAM (.address({address}), .mem_63__7__N_292(mem_63__7__N_292), 
            .data({data}), .mem_60__7__N_283(mem_60__7__N_283), .mem_59__7__N_280(mem_59__7__N_280), 
            .mem_58__7__N_277(mem_58__7__N_277), .mem_56__7__N_271(mem_56__7__N_271), 
            .mem_55__7__N_268(mem_55__7__N_268), .mem_52__7__N_259(mem_52__7__N_259), 
            .mem_51__7__N_256(mem_51__7__N_256), .mem_50__7__N_253(mem_50__7__N_253), 
            .mem_48__7__N_247(mem_48__7__N_247), .mem_47__7__N_244(mem_47__7__N_244), 
            .mem_44__7__N_235(mem_44__7__N_235), .mem_43__7__N_232(mem_43__7__N_232), 
            .mem_42__7__N_229(mem_42__7__N_229), .mem_40__7__N_223(mem_40__7__N_223), 
            .mem_39__7__N_220(mem_39__7__N_220), .mem_36__7__N_211(mem_36__7__N_211), 
            .mem_35__7__N_208(mem_35__7__N_208), .mem_34__7__N_205(mem_34__7__N_205), 
            .mem_32__7__N_199(mem_32__7__N_199), .mem_31__7__N_196(mem_31__7__N_196), 
            .mem_28__7__N_187(mem_28__7__N_187), .mem_27__7__N_184(mem_27__7__N_184), 
            .mem_26__7__N_181(mem_26__7__N_181), .akku_o_c_0(akku_o_c_0), 
            .data_7__N_97(data_7__N_97), .n1905(n1905), .mem_24__7__N_175(mem_24__7__N_175), 
            .mem_23__7__N_172(mem_23__7__N_172), .mem_20__7__N_163(mem_20__7__N_163), 
            .mem_19__7__N_160(mem_19__7__N_160), .mem_18__7__N_157(mem_18__7__N_157), 
            .mem_16__7__N_151(mem_16__7__N_151), .mem_15__7__N_148(mem_15__7__N_148), 
            .mem_12__7__N_139(mem_12__7__N_139), .mem_11__7__N_136(mem_11__7__N_136), 
            .mem_10__7__N_133(mem_10__7__N_133), .mem_8__7__N_127(mem_8__7__N_127), 
            .mem_7__7__N_124(mem_7__7__N_124), .mem_4__7__N_115(mem_4__7__N_115), 
            .mem_3__7__N_112(mem_3__7__N_112), .mem_2__7__N_109(mem_2__7__N_109), 
            .mem_0__7__N_101(mem_0__7__N_101), .akku_o_c_8(akku_o_c_8), 
            .n1895(n1895), .\states_2__N_71[2] (states_2__N_71[2]), .\states_2__N_71[0] (states_2__N_71[0]), 
            .n1302(n1302), .n1898(n1898), .n1896(n1896), .n1906(n1906), 
            .n1902(n1902), .n1901(n1901), .n1911(n1911), .n1910(n1910), 
            .n1899(n1899), .n1900(n1900), .n1327(n1327), .n1328(n1328), 
            .akku_o_c_1(akku_o_c_1), .akku_o_c_2(akku_o_c_2), .akku_o_c_3(akku_o_c_3), 
            .akku_o_c_4(akku_o_c_4), .akku_o_c_5(akku_o_c_5), .akku_o_c_6(akku_o_c_6), 
            .akku_o_c_7(akku_o_c_7), .n1916(n1916));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(44[10:19])
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    CPU8BIT2 CPU (.address({address}), .clk_c(clk_c), .akku_o_c_0(akku_o_c_0), 
            .n1916(n1916), .data({data}), .akku_o_c_7(akku_o_c_7), .akku_o_c_6(akku_o_c_6), 
            .akku_o_c_5(akku_o_c_5), .akku_o_c_4(akku_o_c_4), .\states_2__N_71[2] (states_2__N_71[2]), 
            .akku_o_c_3(akku_o_c_3), .akku_o_c_2(akku_o_c_2), .akku_o_c_1(akku_o_c_1), 
            .reset_c(reset_c), .data_7__N_97(data_7__N_97), .n1895(n1895), 
            .n1905(n1905), .n1328(n1328), .n1898(n1898), .mem_0__7__N_101(mem_0__7__N_101), 
            .n1899(n1899), .mem_15__7__N_148(mem_15__7__N_148), .n1302(n1302), 
            .mem_12__7__N_139(mem_12__7__N_139), .mem_7__7__N_124(mem_7__7__N_124), 
            .n1906(n1906), .mem_56__7__N_271(mem_56__7__N_271), .n1327(n1327), 
            .mem_58__7__N_277(mem_58__7__N_277), .mem_59__7__N_280(mem_59__7__N_280), 
            .mem_60__7__N_283(mem_60__7__N_283), .mem_63__7__N_292(mem_63__7__N_292), 
            .n1902(n1902), .mem_48__7__N_247(mem_48__7__N_247), .mem_50__7__N_253(mem_50__7__N_253), 
            .mem_51__7__N_256(mem_51__7__N_256), .mem_52__7__N_259(mem_52__7__N_259), 
            .mem_55__7__N_268(mem_55__7__N_268), .n1901(n1901), .mem_40__7__N_223(mem_40__7__N_223), 
            .mem_42__7__N_229(mem_42__7__N_229), .mem_43__7__N_232(mem_43__7__N_232), 
            .mem_44__7__N_235(mem_44__7__N_235), .mem_47__7__N_244(mem_47__7__N_244), 
            .n1911(n1911), .mem_32__7__N_199(mem_32__7__N_199), .mem_34__7__N_205(mem_34__7__N_205), 
            .mem_35__7__N_208(mem_35__7__N_208), .mem_36__7__N_211(mem_36__7__N_211), 
            .mem_39__7__N_220(mem_39__7__N_220), .n1910(n1910), .mem_24__7__N_175(mem_24__7__N_175), 
            .mem_26__7__N_181(mem_26__7__N_181), .mem_27__7__N_184(mem_27__7__N_184), 
            .akku_o_c_8(akku_o_c_8), .mem_28__7__N_187(mem_28__7__N_187), 
            .\states_2__N_71[0] (states_2__N_71[0]), .n1896(n1896), .mem_31__7__N_196(mem_31__7__N_196), 
            .n1900(n1900), .mem_16__7__N_151(mem_16__7__N_151), .mem_18__7__N_157(mem_18__7__N_157), 
            .mem_19__7__N_160(mem_19__7__N_160), .mem_20__7__N_163(mem_20__7__N_163), 
            .mem_23__7__N_172(mem_23__7__N_172), .mem_8__7__N_127(mem_8__7__N_127), 
            .mem_10__7__N_133(mem_10__7__N_133), .mem_11__7__N_136(mem_11__7__N_136), 
            .mem_4__7__N_115(mem_4__7__N_115), .mem_3__7__N_112(mem_3__7__N_112), 
            .mem_2__7__N_109(mem_2__7__N_109), .GND_net(GND_net));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(43[10:18])
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module \sram64kx8("sram64kx8.dat")(1,13) 
//

module \sram64kx8("sram64kx8.dat")(1,13)  (address, mem_63__7__N_292, data, 
            mem_60__7__N_283, mem_59__7__N_280, mem_58__7__N_277, mem_56__7__N_271, 
            mem_55__7__N_268, mem_52__7__N_259, mem_51__7__N_256, mem_50__7__N_253, 
            mem_48__7__N_247, mem_47__7__N_244, mem_44__7__N_235, mem_43__7__N_232, 
            mem_42__7__N_229, mem_40__7__N_223, mem_39__7__N_220, mem_36__7__N_211, 
            mem_35__7__N_208, mem_34__7__N_205, mem_32__7__N_199, mem_31__7__N_196, 
            mem_28__7__N_187, mem_27__7__N_184, mem_26__7__N_181, akku_o_c_0, 
            data_7__N_97, n1905, mem_24__7__N_175, mem_23__7__N_172, 
            mem_20__7__N_163, mem_19__7__N_160, mem_18__7__N_157, mem_16__7__N_151, 
            mem_15__7__N_148, mem_12__7__N_139, mem_11__7__N_136, mem_10__7__N_133, 
            mem_8__7__N_127, mem_7__7__N_124, mem_4__7__N_115, mem_3__7__N_112, 
            mem_2__7__N_109, mem_0__7__N_101, akku_o_c_8, n1895, \states_2__N_71[2] , 
            \states_2__N_71[0] , n1302, n1898, n1896, n1906, n1902, 
            n1901, n1911, n1910, n1899, n1900, n1327, n1328, akku_o_c_1, 
            akku_o_c_2, akku_o_c_3, akku_o_c_4, akku_o_c_5, akku_o_c_6, 
            akku_o_c_7, n1916);
    input [5:0]address;
    input mem_63__7__N_292;
    output [7:0]data;
    input mem_60__7__N_283;
    input mem_59__7__N_280;
    input mem_58__7__N_277;
    input mem_56__7__N_271;
    input mem_55__7__N_268;
    input mem_52__7__N_259;
    input mem_51__7__N_256;
    input mem_50__7__N_253;
    input mem_48__7__N_247;
    input mem_47__7__N_244;
    input mem_44__7__N_235;
    input mem_43__7__N_232;
    input mem_42__7__N_229;
    input mem_40__7__N_223;
    input mem_39__7__N_220;
    input mem_36__7__N_211;
    input mem_35__7__N_208;
    input mem_34__7__N_205;
    input mem_32__7__N_199;
    input mem_31__7__N_196;
    input mem_28__7__N_187;
    input mem_27__7__N_184;
    input mem_26__7__N_181;
    input akku_o_c_0;
    input data_7__N_97;
    input n1905;
    input mem_24__7__N_175;
    input mem_23__7__N_172;
    input mem_20__7__N_163;
    input mem_19__7__N_160;
    input mem_18__7__N_157;
    input mem_16__7__N_151;
    input mem_15__7__N_148;
    input mem_12__7__N_139;
    input mem_11__7__N_136;
    input mem_10__7__N_133;
    input mem_8__7__N_127;
    input mem_7__7__N_124;
    input mem_4__7__N_115;
    input mem_3__7__N_112;
    input mem_2__7__N_109;
    input mem_0__7__N_101;
    input akku_o_c_8;
    output n1895;
    output \states_2__N_71[2] ;
    output \states_2__N_71[0] ;
    output n1302;
    output n1898;
    input n1896;
    output n1906;
    output n1902;
    output n1901;
    output n1911;
    output n1910;
    output n1899;
    output n1900;
    output n1327;
    output n1328;
    input akku_o_c_1;
    input akku_o_c_2;
    input akku_o_c_3;
    input akku_o_c_4;
    input akku_o_c_5;
    input akku_o_c_6;
    input akku_o_c_7;
    output n1916;
    
    wire mem_63__7__N_292 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_63__7__N_292 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_62__7__N_289 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_62__7__N_289 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_61__7__N_286 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_61__7__N_286 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_60__7__N_283 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_60__7__N_283 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_59__7__N_280 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_59__7__N_280 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_58__7__N_277 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_58__7__N_277 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_57__7__N_274 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_57__7__N_274 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_56__7__N_271 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_56__7__N_271 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_55__7__N_268 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_55__7__N_268 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_54__7__N_265 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_54__7__N_265 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_53__7__N_262 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_53__7__N_262 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_52__7__N_259 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_52__7__N_259 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_51__7__N_256 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_51__7__N_256 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_50__7__N_253 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_50__7__N_253 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_49__7__N_250 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_49__7__N_250 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_48__7__N_247 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_48__7__N_247 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_47__7__N_244 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_47__7__N_244 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_46__7__N_241 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_46__7__N_241 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_45__7__N_238 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_45__7__N_238 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_44__7__N_235 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_44__7__N_235 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_43__7__N_232 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_43__7__N_232 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_42__7__N_229 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_42__7__N_229 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_41__7__N_226 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_41__7__N_226 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_40__7__N_223 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_40__7__N_223 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_39__7__N_220 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_39__7__N_220 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_38__7__N_217 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_38__7__N_217 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_37__7__N_214 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_37__7__N_214 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_36__7__N_211 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_36__7__N_211 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_35__7__N_208 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_35__7__N_208 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_34__7__N_205 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_34__7__N_205 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_33__7__N_202 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_33__7__N_202 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_32__7__N_199 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_32__7__N_199 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_31__7__N_196 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_31__7__N_196 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_30__7__N_193 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_30__7__N_193 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_29__7__N_190 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_29__7__N_190 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_28__7__N_187 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_28__7__N_187 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_27__7__N_184 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_27__7__N_184 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_26__7__N_181 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_26__7__N_181 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_25__7__N_178 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_25__7__N_178 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_24__7__N_175 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_24__7__N_175 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_23__7__N_172 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_23__7__N_172 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_22__7__N_169 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_22__7__N_169 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_21__7__N_166 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_21__7__N_166 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_20__7__N_163 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_20__7__N_163 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_19__7__N_160 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_19__7__N_160 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_18__7__N_157 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_18__7__N_157 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_17__7__N_154 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_17__7__N_154 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_16__7__N_151 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_16__7__N_151 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_15__7__N_148 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_15__7__N_148 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_14__7__N_145 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_14__7__N_145 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_13__7__N_142 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_13__7__N_142 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_12__7__N_139 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_12__7__N_139 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_11__7__N_136 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_11__7__N_136 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_10__7__N_133 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_10__7__N_133 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_9__7__N_130 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_9__7__N_130 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_8__7__N_127 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_8__7__N_127 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_7__7__N_124 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_7__7__N_124 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_6__7__N_121 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_6__7__N_121 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_5__7__N_118 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_5__7__N_118 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_4__7__N_115 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_4__7__N_115 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_3__7__N_112 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_3__7__N_112 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_2__7__N_109 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_2__7__N_109 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_1__7__N_106 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_1__7__N_106 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_0__7__N_101 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_0__7__N_101 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[16] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[17] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1499;
    wire [7:0]\mem[14] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[15] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1436, n1437;
    wire [7:0]\mem[63] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[18] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[19] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1438;
    wire [7:0]\mem[20] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[21] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1439;
    wire [7:0]\mem[22] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[23] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1440;
    wire [7:0]\mem[48] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[49] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1747, n1501, n1502, n1512;
    wire [7:0]\mem[2] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[3] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1492;
    wire [7:0]\mem[50] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[51] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1748;
    wire [7:0]\mem[24] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[25] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1441, n1784, n1785, n1793;
    wire [7:0]\mem[4] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[5] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1493;
    wire [7:0]\mem[26] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[27] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1442;
    wire [7:0]\mem[28] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[29] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1443;
    wire [7:0]\mem[30] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[31] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1444;
    wire [7:0]\mem[52] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[53] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1749;
    wire [7:0]\mem[54] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[55] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1750;
    wire [7:0]\mem[32] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[33] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1646;
    wire [7:0]\mem[6] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[7] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1494;
    wire [7:0]\mem[8] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[9] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1495;
    wire [7:0]\mem[10] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[11] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1496;
    wire [7:0]\mem[34] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[35] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1647;
    wire [7:0]\mem[56] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[57] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1751;
    wire [7:0]\mem[58] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[59] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1752, n1503, n1504, n1513;
    wire [7:0]\mem[60] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[61] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1753;
    wire [7:0]\mem[36] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[37] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1710, n1709;
    wire [7:0]\mem[62] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1754, n1648, n1708;
    wire [7:0]\mem[38] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[39] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1649;
    wire [7:0]\mem[40] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[41] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1650, n1783, n1505, n1506, n1514, n1805, n1806, n1819, 
        n1677, n1678, n1693, n1679, n1680, n1694, n1681, n1682, 
        n1695, n1807, n1808, n1820, n1809, n1810, n1821, n1683, 
        n1684, n1696;
    wire [7:0]\mem[42] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[43] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1651;
    wire [7:0]\mem[44] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[45] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1652;
    wire [7:0]\mem[46] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[47] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1653, n1654, n1655, n1782, n1656, n1657, n1658;
    wire [7:0]data_7__N_84;
    wire [7:0]\mem[13] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[12] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1659;
    wire [7:0]\mem[0] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[1] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n1460, n1461, n1660, n1661, n1462, n1463, n1685, n1686, 
        n1697, n1464, n1465, n1466, n1568, n1467, n1468, n1687, 
        n1688, n1698, n1469, n1470, n1471, n1472, n1689, n1690, 
        n1699, n1473, n1567, n1474, n1691, n1692, n1700, n1475, 
        n1522, n1523, n1538, n1801, n1524, n1525, n1539, n1802, 
        n1803, n1497, n1498, n1510, n1804, n1491, n1526, n1527, 
        n1540, n1528, n1529, n1541, n1530, n1531, n1542, n1811, 
        n1812, n1822, n1718, n1719, n1729, n1532, n1533, n1543, 
        n1534, n1535, n1544, n1781, n1712, n1713, n1726, n1813, 
        n1814, n1823, n1780, n1536, n1537, n1545, n1345, n1815, 
        n1816, n1824, n1581, n1582, n1583, n1612, n1613, n1614, 
        n1344, n1770, n1771, n1786, n1550, n1551, n1552, n1643, 
        n1644, n1645, n1346, n1347, n1357, n1519, n1520, n1521, 
        n1674, n1675, n1676, n1488, n1489, n1490, n1705, n1706, 
        n1707, n1566, n1457, n1458, n1459, n1736, n1737, n1738, 
        n1426, n1427, n1428, n1767, n1768, n1769, n1395, n1396, 
        n1397, n1798, n1799, n1800, n1364, n1365, n1366, n1829, 
        n1830, n1831, n1772, n1773, n1787, n1584, n1585, n1722, 
        n1723, n1350, n1351, n1586, n1587, n1588, n1589, n1590, 
        n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, 
        n1599, n1367, n1368, n1369, n1370, n1371, n1372, n1373, 
        n1774, n1775, n1788, n1374, n1375, n1376, n1377, n1378, 
        n1379, n1380, n1381, n1382, n1615, n1616, n1617, n1618, 
        n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, 
        n1627, n1628, n1629, n1630, n1565, n1776, n1777, n1789, 
        n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, 
        n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, 
        n1739, n1717, n1553, n1554, n1569, n1740, n1741, n1742, 
        n1743, n1744, n1429, n1720, n1721, n1730, n1430, n1431, 
        n1432, n1745, n1746, n1433, n1434, n1435, n1564, n1714, 
        n1715, n1727, n1349, n1904, n1563, n1555, n1556, n1570, 
        n1562, n1561, n1560, n1559, n1343, n1342, n1341, n1336, 
        n1337, n1352, n1340, n787, n1557, n1558, n1571, n1779, 
        n1348, n1358, n1778, n1338, n1339, n1353, n1790, n1354, 
        n1355, n1572, n1573, n1574, n1575, n1711, n1356, n1716, 
        n1728, n1791, n1576, n1500, n1792, n1724, n1725, n1511, 
        n1509, n1508, n1507, n1818, n1817, n1483, n1482, n1481, 
        n1480, n1479, n1478, n1477, n1669, n1476, n1668, n1667, 
        n1666, n1665, n1664, n1663, n1762, n1761, n1662, n1760, 
        n1452, n1451, n1759, n1450, n1449, n1448, n1447, n1758, 
        n1446, n1445, n1757, n1756, n1755, n1421, n1420, n1419, 
        n1418, n1417, n1416, n1415, n1414, n1638, n1637, n1636, 
        n1635, n1634, n1633, n1632, n1631, n1390, n1389, n1388, 
        n1387, n1386, n1385, n1384, n1383, n1607, n1606, n1605, 
        n1604, n1603, n1602, n1601, n1359, n1731, n1600, n1796, 
        n1795, n1828, n1794, n1580, n1579, n1578, n1577, n1827, 
        n1826, n1825, n1549, n1548, n1547, n1546, n1704, n1703, 
        n1702, n1701, n1518, n1517, n1516, n1515, n1487, n1486, 
        n1485, n1484, n1673, n1672, n1671, n1766, n1670, n1765, 
        n1764, n1763, n1456, n1455, n1454, n1453, n1425, n1424, 
        n1423, n1422, n1642, n1641, n1640, n1639, n1394, n1393, 
        n1392, n1391, n1611, n1610, n1735, n1609, n1608, n1734, 
        n1733, n1363, n1362, n1361, n1732, n1360, n1797;
    
    LUT4 i1313_3_lut (.A(\mem[16] [3]), .B(\mem[17] [3]), .C(address[0]), 
         .Z(n1499)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1313_3_lut.init = 16'hcaca;
    LUT4 i1250_3_lut (.A(\mem[14] [5]), .B(\mem[15] [5]), .C(address[0]), 
         .Z(n1436)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1250_3_lut.init = 16'hcaca;
    LUT4 i1251_3_lut (.A(\mem[16] [5]), .B(\mem[17] [5]), .C(address[0]), 
         .Z(n1437)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1251_3_lut.init = 16'hcaca;
    FD1S1A data_7__I_0_i1 (.D(data[0]), .CK(mem_63__7__N_292), .Q(\mem[63] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i1.GSR = "DISABLED";
    LUT4 i1252_3_lut (.A(\mem[18] [5]), .B(\mem[19] [5]), .C(address[0]), 
         .Z(n1438)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1252_3_lut.init = 16'hcaca;
    LUT4 i1253_3_lut (.A(\mem[20] [5]), .B(\mem[21] [5]), .C(address[0]), 
         .Z(n1439)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1253_3_lut.init = 16'hcaca;
    LUT4 i1254_3_lut (.A(\mem[22] [5]), .B(\mem[23] [5]), .C(address[0]), 
         .Z(n1440)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1254_3_lut.init = 16'hcaca;
    LUT4 i1561_3_lut (.A(\mem[48] [6]), .B(\mem[49] [6]), .C(address[0]), 
         .Z(n1747)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1561_3_lut.init = 16'hcaca;
    PFUMX i1326 (.BLUT(n1501), .ALUT(n1502), .C0(address[1]), .Z(n1512));
    LUT4 i1306_3_lut (.A(\mem[2] [3]), .B(\mem[3] [3]), .C(address[0]), 
         .Z(n1492)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1306_3_lut.init = 16'hcaca;
    LUT4 i1562_3_lut (.A(\mem[50] [6]), .B(\mem[51] [6]), .C(address[0]), 
         .Z(n1748)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1562_3_lut.init = 16'hcaca;
    LUT4 i1255_3_lut (.A(\mem[24] [5]), .B(\mem[25] [5]), .C(address[0]), 
         .Z(n1441)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1255_3_lut.init = 16'hcaca;
    PFUMX i1607 (.BLUT(n1784), .ALUT(n1785), .C0(address[1]), .Z(n1793));
    LUT4 i1307_3_lut (.A(\mem[4] [3]), .B(\mem[5] [3]), .C(address[0]), 
         .Z(n1493)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1307_3_lut.init = 16'hcaca;
    LUT4 i1256_3_lut (.A(\mem[26] [5]), .B(\mem[27] [5]), .C(address[0]), 
         .Z(n1442)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1256_3_lut.init = 16'hcaca;
    LUT4 i1257_3_lut (.A(\mem[28] [5]), .B(\mem[29] [5]), .C(address[0]), 
         .Z(n1443)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1257_3_lut.init = 16'hcaca;
    LUT4 i1258_3_lut (.A(\mem[30] [5]), .B(\mem[31] [5]), .C(address[0]), 
         .Z(n1444)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1258_3_lut.init = 16'hcaca;
    LUT4 i1563_3_lut (.A(\mem[52] [6]), .B(\mem[53] [6]), .C(address[0]), 
         .Z(n1749)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1563_3_lut.init = 16'hcaca;
    LUT4 i1564_3_lut (.A(\mem[54] [6]), .B(\mem[55] [6]), .C(address[0]), 
         .Z(n1750)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1564_3_lut.init = 16'hcaca;
    LUT4 i1460_3_lut (.A(\mem[32] [3]), .B(\mem[33] [3]), .C(address[0]), 
         .Z(n1646)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1460_3_lut.init = 16'hcaca;
    LUT4 i1308_3_lut (.A(\mem[6] [3]), .B(\mem[7] [3]), .C(address[0]), 
         .Z(n1494)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1308_3_lut.init = 16'hcaca;
    LUT4 i1309_3_lut (.A(\mem[8] [3]), .B(\mem[9] [3]), .C(address[0]), 
         .Z(n1495)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1309_3_lut.init = 16'hcaca;
    LUT4 i1310_3_lut (.A(\mem[10] [3]), .B(\mem[11] [3]), .C(address[0]), 
         .Z(n1496)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1310_3_lut.init = 16'hcaca;
    LUT4 i1461_3_lut (.A(\mem[34] [3]), .B(\mem[35] [3]), .C(address[0]), 
         .Z(n1647)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1461_3_lut.init = 16'hcaca;
    LUT4 i1565_3_lut (.A(\mem[56] [6]), .B(\mem[57] [6]), .C(address[0]), 
         .Z(n1751)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1565_3_lut.init = 16'hcaca;
    LUT4 i1566_3_lut (.A(\mem[58] [6]), .B(\mem[59] [6]), .C(address[0]), 
         .Z(n1752)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1566_3_lut.init = 16'hcaca;
    PFUMX i1327 (.BLUT(n1503), .ALUT(n1504), .C0(address[1]), .Z(n1513));
    LUT4 i1567_3_lut (.A(\mem[60] [6]), .B(\mem[61] [6]), .C(address[0]), 
         .Z(n1753)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1567_3_lut.init = 16'hcaca;
    LUT4 i1524_3_lut (.A(\mem[36] [5]), .B(\mem[37] [5]), .C(address[0]), 
         .Z(n1710)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1524_3_lut.init = 16'hcaca;
    LUT4 i1523_3_lut (.A(\mem[34] [5]), .B(\mem[35] [5]), .C(address[0]), 
         .Z(n1709)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1523_3_lut.init = 16'hcaca;
    FD1S1A data_7__I_0_5187_i1 (.D(data[0]), .CK(mem_62__7__N_289), .Q(\mem[62] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i1.GSR = "DISABLED";
    LUT4 i1568_3_lut (.A(\mem[62] [6]), .B(\mem[63] [6]), .C(address[0]), 
         .Z(n1754)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1568_3_lut.init = 16'hcaca;
    LUT4 i1462_3_lut (.A(\mem[36] [3]), .B(\mem[37] [3]), .C(address[0]), 
         .Z(n1648)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1462_3_lut.init = 16'hcaca;
    LUT4 i1522_3_lut (.A(\mem[32] [5]), .B(\mem[33] [5]), .C(address[0]), 
         .Z(n1708)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1522_3_lut.init = 16'hcaca;
    LUT4 i1463_3_lut (.A(\mem[38] [3]), .B(\mem[39] [3]), .C(address[0]), 
         .Z(n1649)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1463_3_lut.init = 16'hcaca;
    LUT4 i1464_3_lut (.A(\mem[40] [3]), .B(\mem[41] [3]), .C(address[0]), 
         .Z(n1650)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1464_3_lut.init = 16'hcaca;
    LUT4 i1597_3_lut (.A(\mem[58] [2]), .B(\mem[59] [2]), .C(address[0]), 
         .Z(n1783)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1597_3_lut.init = 16'hcaca;
    PFUMX i1328 (.BLUT(n1505), .ALUT(n1506), .C0(address[1]), .Z(n1514));
    PFUMX i1633 (.BLUT(n1805), .ALUT(n1806), .C0(address[1]), .Z(n1819));
    PFUMX i1507 (.BLUT(n1677), .ALUT(n1678), .C0(address[1]), .Z(n1693));
    PFUMX i1508 (.BLUT(n1679), .ALUT(n1680), .C0(address[1]), .Z(n1694));
    PFUMX i1509 (.BLUT(n1681), .ALUT(n1682), .C0(address[1]), .Z(n1695));
    PFUMX i1634 (.BLUT(n1807), .ALUT(n1808), .C0(address[1]), .Z(n1820));
    PFUMX i1635 (.BLUT(n1809), .ALUT(n1810), .C0(address[1]), .Z(n1821));
    PFUMX i1510 (.BLUT(n1683), .ALUT(n1684), .C0(address[1]), .Z(n1696));
    LUT4 i1465_3_lut (.A(\mem[42] [3]), .B(\mem[43] [3]), .C(address[0]), 
         .Z(n1651)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1465_3_lut.init = 16'hcaca;
    LUT4 i1466_3_lut (.A(\mem[44] [3]), .B(\mem[45] [3]), .C(address[0]), 
         .Z(n1652)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1466_3_lut.init = 16'hcaca;
    LUT4 i1467_3_lut (.A(\mem[46] [3]), .B(\mem[47] [3]), .C(address[0]), 
         .Z(n1653)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1467_3_lut.init = 16'hcaca;
    LUT4 i1468_3_lut (.A(\mem[48] [3]), .B(\mem[49] [3]), .C(address[0]), 
         .Z(n1654)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1468_3_lut.init = 16'hcaca;
    LUT4 i1469_3_lut (.A(\mem[50] [3]), .B(\mem[51] [3]), .C(address[0]), 
         .Z(n1655)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1469_3_lut.init = 16'hcaca;
    LUT4 i1596_3_lut (.A(\mem[56] [2]), .B(\mem[57] [2]), .C(address[0]), 
         .Z(n1782)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1596_3_lut.init = 16'hcaca;
    LUT4 i1470_3_lut (.A(\mem[52] [3]), .B(\mem[53] [3]), .C(address[0]), 
         .Z(n1656)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1470_3_lut.init = 16'hcaca;
    LUT4 i1471_3_lut (.A(\mem[54] [3]), .B(\mem[55] [3]), .C(address[0]), 
         .Z(n1657)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1471_3_lut.init = 16'hcaca;
    LUT4 i1472_3_lut (.A(\mem[56] [3]), .B(\mem[57] [3]), .C(address[0]), 
         .Z(n1658)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1472_3_lut.init = 16'hcaca;
    FD1S1A data_7__I_0_5184_i1 (.D(data[0]), .CK(mem_61__7__N_286), .Q(\mem[61] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i1 (.D(data[0]), .CK(mem_60__7__N_283), .Q(\mem[60] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i1 (.D(data[0]), .CK(mem_59__7__N_280), .Q(\mem[59] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i1 (.D(data[0]), .CK(mem_58__7__N_277), .Q(\mem[58] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i1 (.D(data[0]), .CK(mem_57__7__N_274), .Q(\mem[57] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i1 (.D(data[0]), .CK(mem_56__7__N_271), .Q(\mem[56] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i1 (.D(data[0]), .CK(mem_55__7__N_268), .Q(\mem[55] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i1 (.D(data[0]), .CK(mem_54__7__N_265), .Q(\mem[54] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i1 (.D(data[0]), .CK(mem_53__7__N_262), .Q(\mem[53] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i1 (.D(data[0]), .CK(mem_52__7__N_259), .Q(\mem[52] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i1 (.D(data[0]), .CK(mem_51__7__N_256), .Q(\mem[51] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i1 (.D(data[0]), .CK(mem_50__7__N_253), .Q(\mem[50] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i1 (.D(data[0]), .CK(mem_49__7__N_250), .Q(\mem[49] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i1 (.D(data[0]), .CK(mem_48__7__N_247), .Q(\mem[48] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i1 (.D(data[0]), .CK(mem_47__7__N_244), .Q(\mem[47] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i1 (.D(data[0]), .CK(mem_46__7__N_241), .Q(\mem[46] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i1 (.D(data[0]), .CK(mem_45__7__N_238), .Q(\mem[45] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i1 (.D(data[0]), .CK(mem_44__7__N_235), .Q(\mem[44] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i1 (.D(data[0]), .CK(mem_43__7__N_232), .Q(\mem[43] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i1 (.D(data[0]), .CK(mem_42__7__N_229), .Q(\mem[42] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i1 (.D(data[0]), .CK(mem_41__7__N_226), .Q(\mem[41] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i1 (.D(data[0]), .CK(mem_40__7__N_223), .Q(\mem[40] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i1 (.D(data[0]), .CK(mem_39__7__N_220), .Q(\mem[39] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i1 (.D(data[0]), .CK(mem_38__7__N_217), .Q(\mem[38] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i1 (.D(data[0]), .CK(mem_37__7__N_214), .Q(\mem[37] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i1 (.D(data[0]), .CK(mem_36__7__N_211), .Q(\mem[36] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i1 (.D(data[0]), .CK(mem_35__7__N_208), .Q(\mem[35] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i1 (.D(data[0]), .CK(mem_34__7__N_205), .Q(\mem[34] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i1 (.D(data[0]), .CK(mem_33__7__N_202), .Q(\mem[33] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i1 (.D(data[0]), .CK(mem_32__7__N_199), .Q(\mem[32] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i1 (.D(data[0]), .CK(mem_31__7__N_196), .Q(\mem[31] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i1 (.D(data[0]), .CK(mem_30__7__N_193), .Q(\mem[30] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i1 (.D(data[0]), .CK(mem_29__7__N_190), .Q(\mem[29] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i1 (.D(data[0]), .CK(mem_28__7__N_187), .Q(\mem[28] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i1 (.D(data[0]), .CK(mem_27__7__N_184), .Q(\mem[27] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i1 (.D(data[0]), .CK(mem_26__7__N_181), .Q(\mem[26] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i1 (.D(data[0]), .CK(mem_25__7__N_178), .Q(\mem[25] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i1.GSR = "DISABLED";
    LUT4 Select_407_i3_4_lut (.A(data_7__N_84[0]), .B(akku_o_c_0), .C(data_7__N_97), 
         .D(n1905), .Z(data[0])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_407_i3_4_lut.init = 16'ha0ec;
    FD1S1A data_7__I_0_5073_i1 (.D(data[0]), .CK(mem_24__7__N_175), .Q(\mem[24] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i1 (.D(data[0]), .CK(mem_23__7__N_172), .Q(\mem[23] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i1 (.D(data[0]), .CK(mem_22__7__N_169), .Q(\mem[22] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i1 (.D(data[0]), .CK(mem_21__7__N_166), .Q(\mem[21] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5061_i1 (.D(data[0]), .CK(mem_20__7__N_163), .Q(\mem[20] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i1 (.D(data[0]), .CK(mem_19__7__N_160), .Q(\mem[19] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5055_i1 (.D(data[0]), .CK(mem_18__7__N_157), .Q(\mem[18] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5052_i1 (.D(data[0]), .CK(mem_17__7__N_154), .Q(\mem[17] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i1 (.D(data[0]), .CK(mem_16__7__N_151), .Q(\mem[16] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5046_i1 (.D(data[0]), .CK(mem_15__7__N_148), .Q(\mem[15] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5043_i1 (.D(data[0]), .CK(mem_14__7__N_145), .Q(\mem[14] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5040_i1 (.D(data[0]), .CK(mem_13__7__N_142), .Q(\mem[13] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5037_i1 (.D(data[0]), .CK(mem_12__7__N_139), .Q(\mem[12] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i1 (.D(data[0]), .CK(mem_11__7__N_136), .Q(\mem[11] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i1.GSR = "DISABLED";
    LUT4 i1473_3_lut (.A(\mem[58] [3]), .B(\mem[59] [3]), .C(address[0]), 
         .Z(n1659)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1473_3_lut.init = 16'hcaca;
    LUT4 i1274_3_lut (.A(\mem[0] [4]), .B(\mem[1] [4]), .C(address[0]), 
         .Z(n1460)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1274_3_lut.init = 16'hcaca;
    FD1S1A data_7__I_0_5031_i1 (.D(data[0]), .CK(mem_10__7__N_133), .Q(\mem[10] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5028_i1 (.D(data[0]), .CK(mem_9__7__N_130), .Q(\mem[9] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5025_i1 (.D(data[0]), .CK(mem_8__7__N_127), .Q(\mem[8] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5022_i1 (.D(data[0]), .CK(mem_7__7__N_124), .Q(\mem[7] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5019_i1 (.D(data[0]), .CK(mem_6__7__N_121), .Q(\mem[6] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5016_i1 (.D(data[0]), .CK(mem_5__7__N_118), .Q(\mem[5] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5013_i1 (.D(data[0]), .CK(mem_4__7__N_115), .Q(\mem[4] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i1.GSR = "DISABLED";
    LUT4 i1275_3_lut (.A(\mem[2] [4]), .B(\mem[3] [4]), .C(address[0]), 
         .Z(n1461)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1275_3_lut.init = 16'hcaca;
    FD1S1AY data_7__I_0_5010_i1 (.D(data[0]), .CK(mem_3__7__N_112), .Q(\mem[3] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i1.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5007_i1 (.D(data[0]), .CK(mem_2__7__N_109), .Q(\mem[2] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5004_i1 (.D(data[0]), .CK(mem_1__7__N_106), .Q(\mem[1] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i1.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5002_i1 (.D(data[0]), .CK(mem_0__7__N_101), .Q(\mem[0] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i1.GSR = "DISABLED";
    LUT4 i1474_3_lut (.A(\mem[60] [3]), .B(\mem[61] [3]), .C(address[0]), 
         .Z(n1660)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1474_3_lut.init = 16'hcaca;
    LUT4 i1475_3_lut (.A(\mem[62] [3]), .B(\mem[63] [3]), .C(address[0]), 
         .Z(n1661)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1475_3_lut.init = 16'hcaca;
    FD1S1AY data_7__I_0_5002_i2 (.D(data[1]), .CK(mem_0__7__N_101), .Q(\mem[0] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5002_i3 (.D(data[2]), .CK(mem_0__7__N_101), .Q(\mem[0] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5002_i4 (.D(data[3]), .CK(mem_0__7__N_101), .Q(\mem[0] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i4.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5002_i5 (.D(data[4]), .CK(mem_0__7__N_101), .Q(\mem[0] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i5.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5002_i6 (.D(data[5]), .CK(mem_0__7__N_101), .Q(\mem[0] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5002_i7 (.D(data[6]), .CK(mem_0__7__N_101), .Q(\mem[0] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i7.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5002_i8 (.D(data[7]), .CK(mem_0__7__N_101), .Q(\mem[0] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i8.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5004_i2 (.D(data[1]), .CK(mem_1__7__N_106), .Q(\mem[1] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5004_i3 (.D(data[2]), .CK(mem_1__7__N_106), .Q(\mem[1] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5004_i4 (.D(data[3]), .CK(mem_1__7__N_106), .Q(\mem[1] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5004_i5 (.D(data[4]), .CK(mem_1__7__N_106), .Q(\mem[1] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i5.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5004_i6 (.D(data[5]), .CK(mem_1__7__N_106), .Q(\mem[1] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i6.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5004_i7 (.D(data[6]), .CK(mem_1__7__N_106), .Q(\mem[1] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i7.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5004_i8 (.D(data[7]), .CK(mem_1__7__N_106), .Q(\mem[1] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i8.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5007_i2 (.D(data[1]), .CK(mem_2__7__N_109), .Q(\mem[2] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5007_i3 (.D(data[2]), .CK(mem_2__7__N_109), .Q(\mem[2] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i3.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5007_i4 (.D(data[3]), .CK(mem_2__7__N_109), .Q(\mem[2] [3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i4.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5007_i5 (.D(data[4]), .CK(mem_2__7__N_109), .Q(\mem[2] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i5.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5007_i6 (.D(data[5]), .CK(mem_2__7__N_109), .Q(\mem[2] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5007_i7 (.D(data[6]), .CK(mem_2__7__N_109), .Q(\mem[2] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i7.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5007_i8 (.D(data[7]), .CK(mem_2__7__N_109), .Q(\mem[2] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5010_i2 (.D(data[1]), .CK(mem_3__7__N_112), .Q(\mem[3] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5010_i3 (.D(data[2]), .CK(mem_3__7__N_112), .Q(\mem[3] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5010_i4 (.D(data[3]), .CK(mem_3__7__N_112), .Q(\mem[3] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i4.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5010_i5 (.D(data[4]), .CK(mem_3__7__N_112), .Q(\mem[3] [4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i5.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5010_i6 (.D(data[5]), .CK(mem_3__7__N_112), .Q(\mem[3] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i6.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5010_i7 (.D(data[6]), .CK(mem_3__7__N_112), .Q(\mem[3] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i7.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5010_i8 (.D(data[7]), .CK(mem_3__7__N_112), .Q(\mem[3] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5013_i2 (.D(data[1]), .CK(mem_4__7__N_115), .Q(\mem[4] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5013_i3 (.D(data[2]), .CK(mem_4__7__N_115), .Q(\mem[4] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5013_i4 (.D(data[3]), .CK(mem_4__7__N_115), .Q(\mem[4] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5013_i5 (.D(data[4]), .CK(mem_4__7__N_115), .Q(\mem[4] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5013_i6 (.D(data[5]), .CK(mem_4__7__N_115), .Q(\mem[4] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i6.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5013_i7 (.D(data[6]), .CK(mem_4__7__N_115), .Q(\mem[4] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i7.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5013_i8 (.D(data[7]), .CK(mem_4__7__N_115), .Q(\mem[4] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i8.GSR = "DISABLED";
    LUT4 i1276_3_lut (.A(\mem[4] [4]), .B(\mem[5] [4]), .C(address[0]), 
         .Z(n1462)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1276_3_lut.init = 16'hcaca;
    FD1S1A data_7__I_0_i2 (.D(data[1]), .CK(mem_63__7__N_292), .Q(\mem[63] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i2.GSR = "DISABLED";
    LUT4 i1277_3_lut (.A(\mem[6] [4]), .B(\mem[7] [4]), .C(address[0]), 
         .Z(n1463)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1277_3_lut.init = 16'hcaca;
    PFUMX i1511 (.BLUT(n1685), .ALUT(n1686), .C0(address[1]), .Z(n1697));
    FD1S1A data_7__I_0_i3 (.D(data[2]), .CK(mem_63__7__N_292), .Q(\mem[63] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_i4 (.D(data[3]), .CK(mem_63__7__N_292), .Q(\mem[63] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_i5 (.D(data[4]), .CK(mem_63__7__N_292), .Q(\mem[63] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_i6 (.D(data[5]), .CK(mem_63__7__N_292), .Q(\mem[63] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_i7 (.D(data[6]), .CK(mem_63__7__N_292), .Q(\mem[63] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_i8 (.D(data[7]), .CK(mem_63__7__N_292), .Q(\mem[63] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5187_i2 (.D(data[1]), .CK(mem_62__7__N_289), .Q(\mem[62] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5187_i3 (.D(data[2]), .CK(mem_62__7__N_289), .Q(\mem[62] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5187_i4 (.D(data[3]), .CK(mem_62__7__N_289), .Q(\mem[62] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5187_i5 (.D(data[4]), .CK(mem_62__7__N_289), .Q(\mem[62] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5187_i6 (.D(data[5]), .CK(mem_62__7__N_289), .Q(\mem[62] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5187_i7 (.D(data[6]), .CK(mem_62__7__N_289), .Q(\mem[62] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5187_i8 (.D(data[7]), .CK(mem_62__7__N_289), .Q(\mem[62] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i2 (.D(data[1]), .CK(mem_61__7__N_286), .Q(\mem[61] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i3 (.D(data[2]), .CK(mem_61__7__N_286), .Q(\mem[61] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i4 (.D(data[3]), .CK(mem_61__7__N_286), .Q(\mem[61] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i5 (.D(data[4]), .CK(mem_61__7__N_286), .Q(\mem[61] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i6 (.D(data[5]), .CK(mem_61__7__N_286), .Q(\mem[61] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i7 (.D(data[6]), .CK(mem_61__7__N_286), .Q(\mem[61] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i8 (.D(data[7]), .CK(mem_61__7__N_286), .Q(\mem[61] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i2 (.D(data[1]), .CK(mem_60__7__N_283), .Q(\mem[60] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i3 (.D(data[2]), .CK(mem_60__7__N_283), .Q(\mem[60] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i4 (.D(data[3]), .CK(mem_60__7__N_283), .Q(\mem[60] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i5 (.D(data[4]), .CK(mem_60__7__N_283), .Q(\mem[60] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i6 (.D(data[5]), .CK(mem_60__7__N_283), .Q(\mem[60] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i7 (.D(data[6]), .CK(mem_60__7__N_283), .Q(\mem[60] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i8 (.D(data[7]), .CK(mem_60__7__N_283), .Q(\mem[60] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i2 (.D(data[1]), .CK(mem_59__7__N_280), .Q(\mem[59] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i3 (.D(data[2]), .CK(mem_59__7__N_280), .Q(\mem[59] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i4 (.D(data[3]), .CK(mem_59__7__N_280), .Q(\mem[59] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i5 (.D(data[4]), .CK(mem_59__7__N_280), .Q(\mem[59] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i6 (.D(data[5]), .CK(mem_59__7__N_280), .Q(\mem[59] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i7 (.D(data[6]), .CK(mem_59__7__N_280), .Q(\mem[59] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i8 (.D(data[7]), .CK(mem_59__7__N_280), .Q(\mem[59] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i2 (.D(data[1]), .CK(mem_58__7__N_277), .Q(\mem[58] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i3 (.D(data[2]), .CK(mem_58__7__N_277), .Q(\mem[58] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i4 (.D(data[3]), .CK(mem_58__7__N_277), .Q(\mem[58] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i5 (.D(data[4]), .CK(mem_58__7__N_277), .Q(\mem[58] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i6 (.D(data[5]), .CK(mem_58__7__N_277), .Q(\mem[58] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i7 (.D(data[6]), .CK(mem_58__7__N_277), .Q(\mem[58] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i8 (.D(data[7]), .CK(mem_58__7__N_277), .Q(\mem[58] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i2 (.D(data[1]), .CK(mem_57__7__N_274), .Q(\mem[57] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i3 (.D(data[2]), .CK(mem_57__7__N_274), .Q(\mem[57] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i4 (.D(data[3]), .CK(mem_57__7__N_274), .Q(\mem[57] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i5 (.D(data[4]), .CK(mem_57__7__N_274), .Q(\mem[57] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i6 (.D(data[5]), .CK(mem_57__7__N_274), .Q(\mem[57] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i7 (.D(data[6]), .CK(mem_57__7__N_274), .Q(\mem[57] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i8 (.D(data[7]), .CK(mem_57__7__N_274), .Q(\mem[57] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i2 (.D(data[1]), .CK(mem_56__7__N_271), .Q(\mem[56] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i3 (.D(data[2]), .CK(mem_56__7__N_271), .Q(\mem[56] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i4 (.D(data[3]), .CK(mem_56__7__N_271), .Q(\mem[56] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i5 (.D(data[4]), .CK(mem_56__7__N_271), .Q(\mem[56] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i6 (.D(data[5]), .CK(mem_56__7__N_271), .Q(\mem[56] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i7 (.D(data[6]), .CK(mem_56__7__N_271), .Q(\mem[56] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i8 (.D(data[7]), .CK(mem_56__7__N_271), .Q(\mem[56] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i2 (.D(data[1]), .CK(mem_55__7__N_268), .Q(\mem[55] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i3 (.D(data[2]), .CK(mem_55__7__N_268), .Q(\mem[55] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i4 (.D(data[3]), .CK(mem_55__7__N_268), .Q(\mem[55] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i5 (.D(data[4]), .CK(mem_55__7__N_268), .Q(\mem[55] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i6 (.D(data[5]), .CK(mem_55__7__N_268), .Q(\mem[55] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i7 (.D(data[6]), .CK(mem_55__7__N_268), .Q(\mem[55] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i8 (.D(data[7]), .CK(mem_55__7__N_268), .Q(\mem[55] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i2 (.D(data[1]), .CK(mem_54__7__N_265), .Q(\mem[54] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i3 (.D(data[2]), .CK(mem_54__7__N_265), .Q(\mem[54] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i4 (.D(data[3]), .CK(mem_54__7__N_265), .Q(\mem[54] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i5 (.D(data[4]), .CK(mem_54__7__N_265), .Q(\mem[54] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i6 (.D(data[5]), .CK(mem_54__7__N_265), .Q(\mem[54] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i7 (.D(data[6]), .CK(mem_54__7__N_265), .Q(\mem[54] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i8 (.D(data[7]), .CK(mem_54__7__N_265), .Q(\mem[54] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i2 (.D(data[1]), .CK(mem_53__7__N_262), .Q(\mem[53] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i3 (.D(data[2]), .CK(mem_53__7__N_262), .Q(\mem[53] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i4 (.D(data[3]), .CK(mem_53__7__N_262), .Q(\mem[53] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i5 (.D(data[4]), .CK(mem_53__7__N_262), .Q(\mem[53] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i6 (.D(data[5]), .CK(mem_53__7__N_262), .Q(\mem[53] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i7 (.D(data[6]), .CK(mem_53__7__N_262), .Q(\mem[53] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i8 (.D(data[7]), .CK(mem_53__7__N_262), .Q(\mem[53] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i2 (.D(data[1]), .CK(mem_52__7__N_259), .Q(\mem[52] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i3 (.D(data[2]), .CK(mem_52__7__N_259), .Q(\mem[52] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i4 (.D(data[3]), .CK(mem_52__7__N_259), .Q(\mem[52] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i5 (.D(data[4]), .CK(mem_52__7__N_259), .Q(\mem[52] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i6 (.D(data[5]), .CK(mem_52__7__N_259), .Q(\mem[52] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i7 (.D(data[6]), .CK(mem_52__7__N_259), .Q(\mem[52] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i8 (.D(data[7]), .CK(mem_52__7__N_259), .Q(\mem[52] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i2 (.D(data[1]), .CK(mem_51__7__N_256), .Q(\mem[51] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i3 (.D(data[2]), .CK(mem_51__7__N_256), .Q(\mem[51] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i4 (.D(data[3]), .CK(mem_51__7__N_256), .Q(\mem[51] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i5 (.D(data[4]), .CK(mem_51__7__N_256), .Q(\mem[51] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i6 (.D(data[5]), .CK(mem_51__7__N_256), .Q(\mem[51] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i7 (.D(data[6]), .CK(mem_51__7__N_256), .Q(\mem[51] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i8 (.D(data[7]), .CK(mem_51__7__N_256), .Q(\mem[51] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i2 (.D(data[1]), .CK(mem_50__7__N_253), .Q(\mem[50] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i3 (.D(data[2]), .CK(mem_50__7__N_253), .Q(\mem[50] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i4 (.D(data[3]), .CK(mem_50__7__N_253), .Q(\mem[50] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i5 (.D(data[4]), .CK(mem_50__7__N_253), .Q(\mem[50] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i6 (.D(data[5]), .CK(mem_50__7__N_253), .Q(\mem[50] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i7 (.D(data[6]), .CK(mem_50__7__N_253), .Q(\mem[50] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i8 (.D(data[7]), .CK(mem_50__7__N_253), .Q(\mem[50] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i2 (.D(data[1]), .CK(mem_49__7__N_250), .Q(\mem[49] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i3 (.D(data[2]), .CK(mem_49__7__N_250), .Q(\mem[49] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i4 (.D(data[3]), .CK(mem_49__7__N_250), .Q(\mem[49] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i5 (.D(data[4]), .CK(mem_49__7__N_250), .Q(\mem[49] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i6 (.D(data[5]), .CK(mem_49__7__N_250), .Q(\mem[49] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i7 (.D(data[6]), .CK(mem_49__7__N_250), .Q(\mem[49] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i8 (.D(data[7]), .CK(mem_49__7__N_250), .Q(\mem[49] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i2 (.D(data[1]), .CK(mem_48__7__N_247), .Q(\mem[48] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i3 (.D(data[2]), .CK(mem_48__7__N_247), .Q(\mem[48] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i4 (.D(data[3]), .CK(mem_48__7__N_247), .Q(\mem[48] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i5 (.D(data[4]), .CK(mem_48__7__N_247), .Q(\mem[48] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i6 (.D(data[5]), .CK(mem_48__7__N_247), .Q(\mem[48] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i7 (.D(data[6]), .CK(mem_48__7__N_247), .Q(\mem[48] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i8 (.D(data[7]), .CK(mem_48__7__N_247), .Q(\mem[48] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i2 (.D(data[1]), .CK(mem_47__7__N_244), .Q(\mem[47] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i3 (.D(data[2]), .CK(mem_47__7__N_244), .Q(\mem[47] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i4 (.D(data[3]), .CK(mem_47__7__N_244), .Q(\mem[47] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i5 (.D(data[4]), .CK(mem_47__7__N_244), .Q(\mem[47] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i6 (.D(data[5]), .CK(mem_47__7__N_244), .Q(\mem[47] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i7 (.D(data[6]), .CK(mem_47__7__N_244), .Q(\mem[47] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i8 (.D(data[7]), .CK(mem_47__7__N_244), .Q(\mem[47] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i2 (.D(data[1]), .CK(mem_46__7__N_241), .Q(\mem[46] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i3 (.D(data[2]), .CK(mem_46__7__N_241), .Q(\mem[46] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i4 (.D(data[3]), .CK(mem_46__7__N_241), .Q(\mem[46] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i5 (.D(data[4]), .CK(mem_46__7__N_241), .Q(\mem[46] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i6 (.D(data[5]), .CK(mem_46__7__N_241), .Q(\mem[46] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i7 (.D(data[6]), .CK(mem_46__7__N_241), .Q(\mem[46] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i8 (.D(data[7]), .CK(mem_46__7__N_241), .Q(\mem[46] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i2 (.D(data[1]), .CK(mem_45__7__N_238), .Q(\mem[45] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i3 (.D(data[2]), .CK(mem_45__7__N_238), .Q(\mem[45] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i4 (.D(data[3]), .CK(mem_45__7__N_238), .Q(\mem[45] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i5 (.D(data[4]), .CK(mem_45__7__N_238), .Q(\mem[45] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i6 (.D(data[5]), .CK(mem_45__7__N_238), .Q(\mem[45] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i7 (.D(data[6]), .CK(mem_45__7__N_238), .Q(\mem[45] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i8 (.D(data[7]), .CK(mem_45__7__N_238), .Q(\mem[45] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i2 (.D(data[1]), .CK(mem_44__7__N_235), .Q(\mem[44] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i3 (.D(data[2]), .CK(mem_44__7__N_235), .Q(\mem[44] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i4 (.D(data[3]), .CK(mem_44__7__N_235), .Q(\mem[44] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i5 (.D(data[4]), .CK(mem_44__7__N_235), .Q(\mem[44] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i6 (.D(data[5]), .CK(mem_44__7__N_235), .Q(\mem[44] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i7 (.D(data[6]), .CK(mem_44__7__N_235), .Q(\mem[44] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i8 (.D(data[7]), .CK(mem_44__7__N_235), .Q(\mem[44] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i2 (.D(data[1]), .CK(mem_43__7__N_232), .Q(\mem[43] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i3 (.D(data[2]), .CK(mem_43__7__N_232), .Q(\mem[43] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i4 (.D(data[3]), .CK(mem_43__7__N_232), .Q(\mem[43] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i5 (.D(data[4]), .CK(mem_43__7__N_232), .Q(\mem[43] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i6 (.D(data[5]), .CK(mem_43__7__N_232), .Q(\mem[43] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i7 (.D(data[6]), .CK(mem_43__7__N_232), .Q(\mem[43] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i8 (.D(data[7]), .CK(mem_43__7__N_232), .Q(\mem[43] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i2 (.D(data[1]), .CK(mem_42__7__N_229), .Q(\mem[42] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i3 (.D(data[2]), .CK(mem_42__7__N_229), .Q(\mem[42] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i4 (.D(data[3]), .CK(mem_42__7__N_229), .Q(\mem[42] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i5 (.D(data[4]), .CK(mem_42__7__N_229), .Q(\mem[42] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i6 (.D(data[5]), .CK(mem_42__7__N_229), .Q(\mem[42] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i7 (.D(data[6]), .CK(mem_42__7__N_229), .Q(\mem[42] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i8 (.D(data[7]), .CK(mem_42__7__N_229), .Q(\mem[42] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i2 (.D(data[1]), .CK(mem_41__7__N_226), .Q(\mem[41] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i3 (.D(data[2]), .CK(mem_41__7__N_226), .Q(\mem[41] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i4 (.D(data[3]), .CK(mem_41__7__N_226), .Q(\mem[41] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i5 (.D(data[4]), .CK(mem_41__7__N_226), .Q(\mem[41] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i6 (.D(data[5]), .CK(mem_41__7__N_226), .Q(\mem[41] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i7 (.D(data[6]), .CK(mem_41__7__N_226), .Q(\mem[41] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i8 (.D(data[7]), .CK(mem_41__7__N_226), .Q(\mem[41] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i2 (.D(data[1]), .CK(mem_40__7__N_223), .Q(\mem[40] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i3 (.D(data[2]), .CK(mem_40__7__N_223), .Q(\mem[40] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i4 (.D(data[3]), .CK(mem_40__7__N_223), .Q(\mem[40] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i5 (.D(data[4]), .CK(mem_40__7__N_223), .Q(\mem[40] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i6 (.D(data[5]), .CK(mem_40__7__N_223), .Q(\mem[40] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i7 (.D(data[6]), .CK(mem_40__7__N_223), .Q(\mem[40] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i8 (.D(data[7]), .CK(mem_40__7__N_223), .Q(\mem[40] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i2 (.D(data[1]), .CK(mem_39__7__N_220), .Q(\mem[39] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i3 (.D(data[2]), .CK(mem_39__7__N_220), .Q(\mem[39] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i4 (.D(data[3]), .CK(mem_39__7__N_220), .Q(\mem[39] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i5 (.D(data[4]), .CK(mem_39__7__N_220), .Q(\mem[39] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i6 (.D(data[5]), .CK(mem_39__7__N_220), .Q(\mem[39] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i7 (.D(data[6]), .CK(mem_39__7__N_220), .Q(\mem[39] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i8 (.D(data[7]), .CK(mem_39__7__N_220), .Q(\mem[39] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i2 (.D(data[1]), .CK(mem_38__7__N_217), .Q(\mem[38] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i3 (.D(data[2]), .CK(mem_38__7__N_217), .Q(\mem[38] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i4 (.D(data[3]), .CK(mem_38__7__N_217), .Q(\mem[38] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i5 (.D(data[4]), .CK(mem_38__7__N_217), .Q(\mem[38] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i6 (.D(data[5]), .CK(mem_38__7__N_217), .Q(\mem[38] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i7 (.D(data[6]), .CK(mem_38__7__N_217), .Q(\mem[38] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i8 (.D(data[7]), .CK(mem_38__7__N_217), .Q(\mem[38] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i2 (.D(data[1]), .CK(mem_37__7__N_214), .Q(\mem[37] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i3 (.D(data[2]), .CK(mem_37__7__N_214), .Q(\mem[37] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i4 (.D(data[3]), .CK(mem_37__7__N_214), .Q(\mem[37] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i5 (.D(data[4]), .CK(mem_37__7__N_214), .Q(\mem[37] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i6 (.D(data[5]), .CK(mem_37__7__N_214), .Q(\mem[37] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i7 (.D(data[6]), .CK(mem_37__7__N_214), .Q(\mem[37] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i8 (.D(data[7]), .CK(mem_37__7__N_214), .Q(\mem[37] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i2 (.D(data[1]), .CK(mem_36__7__N_211), .Q(\mem[36] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i3 (.D(data[2]), .CK(mem_36__7__N_211), .Q(\mem[36] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i4 (.D(data[3]), .CK(mem_36__7__N_211), .Q(\mem[36] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i5 (.D(data[4]), .CK(mem_36__7__N_211), .Q(\mem[36] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i6 (.D(data[5]), .CK(mem_36__7__N_211), .Q(\mem[36] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i7 (.D(data[6]), .CK(mem_36__7__N_211), .Q(\mem[36] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i8 (.D(data[7]), .CK(mem_36__7__N_211), .Q(\mem[36] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i2 (.D(data[1]), .CK(mem_35__7__N_208), .Q(\mem[35] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i3 (.D(data[2]), .CK(mem_35__7__N_208), .Q(\mem[35] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i4 (.D(data[3]), .CK(mem_35__7__N_208), .Q(\mem[35] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i5 (.D(data[4]), .CK(mem_35__7__N_208), .Q(\mem[35] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i6 (.D(data[5]), .CK(mem_35__7__N_208), .Q(\mem[35] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i7 (.D(data[6]), .CK(mem_35__7__N_208), .Q(\mem[35] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i8 (.D(data[7]), .CK(mem_35__7__N_208), .Q(\mem[35] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i2 (.D(data[1]), .CK(mem_34__7__N_205), .Q(\mem[34] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i3 (.D(data[2]), .CK(mem_34__7__N_205), .Q(\mem[34] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i4 (.D(data[3]), .CK(mem_34__7__N_205), .Q(\mem[34] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i5 (.D(data[4]), .CK(mem_34__7__N_205), .Q(\mem[34] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i6 (.D(data[5]), .CK(mem_34__7__N_205), .Q(\mem[34] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i7 (.D(data[6]), .CK(mem_34__7__N_205), .Q(\mem[34] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i8 (.D(data[7]), .CK(mem_34__7__N_205), .Q(\mem[34] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i2 (.D(data[1]), .CK(mem_33__7__N_202), .Q(\mem[33] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i3 (.D(data[2]), .CK(mem_33__7__N_202), .Q(\mem[33] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i4 (.D(data[3]), .CK(mem_33__7__N_202), .Q(\mem[33] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i5 (.D(data[4]), .CK(mem_33__7__N_202), .Q(\mem[33] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i6 (.D(data[5]), .CK(mem_33__7__N_202), .Q(\mem[33] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i7 (.D(data[6]), .CK(mem_33__7__N_202), .Q(\mem[33] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i8 (.D(data[7]), .CK(mem_33__7__N_202), .Q(\mem[33] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i2 (.D(data[1]), .CK(mem_32__7__N_199), .Q(\mem[32] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i3 (.D(data[2]), .CK(mem_32__7__N_199), .Q(\mem[32] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i4 (.D(data[3]), .CK(mem_32__7__N_199), .Q(\mem[32] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i5 (.D(data[4]), .CK(mem_32__7__N_199), .Q(\mem[32] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i6 (.D(data[5]), .CK(mem_32__7__N_199), .Q(\mem[32] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i7 (.D(data[6]), .CK(mem_32__7__N_199), .Q(\mem[32] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i8 (.D(data[7]), .CK(mem_32__7__N_199), .Q(\mem[32] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i2 (.D(data[1]), .CK(mem_31__7__N_196), .Q(\mem[31] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i3 (.D(data[2]), .CK(mem_31__7__N_196), .Q(\mem[31] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i4 (.D(data[3]), .CK(mem_31__7__N_196), .Q(\mem[31] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i5 (.D(data[4]), .CK(mem_31__7__N_196), .Q(\mem[31] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i6 (.D(data[5]), .CK(mem_31__7__N_196), .Q(\mem[31] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i7 (.D(data[6]), .CK(mem_31__7__N_196), .Q(\mem[31] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i8 (.D(data[7]), .CK(mem_31__7__N_196), .Q(\mem[31] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i2 (.D(data[1]), .CK(mem_30__7__N_193), .Q(\mem[30] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i3 (.D(data[2]), .CK(mem_30__7__N_193), .Q(\mem[30] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i4 (.D(data[3]), .CK(mem_30__7__N_193), .Q(\mem[30] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i5 (.D(data[4]), .CK(mem_30__7__N_193), .Q(\mem[30] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i6 (.D(data[5]), .CK(mem_30__7__N_193), .Q(\mem[30] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i7 (.D(data[6]), .CK(mem_30__7__N_193), .Q(\mem[30] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i8 (.D(data[7]), .CK(mem_30__7__N_193), .Q(\mem[30] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i2 (.D(data[1]), .CK(mem_29__7__N_190), .Q(\mem[29] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i3 (.D(data[2]), .CK(mem_29__7__N_190), .Q(\mem[29] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i4 (.D(data[3]), .CK(mem_29__7__N_190), .Q(\mem[29] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i5 (.D(data[4]), .CK(mem_29__7__N_190), .Q(\mem[29] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i6 (.D(data[5]), .CK(mem_29__7__N_190), .Q(\mem[29] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i7 (.D(data[6]), .CK(mem_29__7__N_190), .Q(\mem[29] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i8 (.D(data[7]), .CK(mem_29__7__N_190), .Q(\mem[29] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i2 (.D(data[1]), .CK(mem_28__7__N_187), .Q(\mem[28] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i3 (.D(data[2]), .CK(mem_28__7__N_187), .Q(\mem[28] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i4 (.D(data[3]), .CK(mem_28__7__N_187), .Q(\mem[28] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i5 (.D(data[4]), .CK(mem_28__7__N_187), .Q(\mem[28] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i6 (.D(data[5]), .CK(mem_28__7__N_187), .Q(\mem[28] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i7 (.D(data[6]), .CK(mem_28__7__N_187), .Q(\mem[28] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i8 (.D(data[7]), .CK(mem_28__7__N_187), .Q(\mem[28] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i2 (.D(data[1]), .CK(mem_27__7__N_184), .Q(\mem[27] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i3 (.D(data[2]), .CK(mem_27__7__N_184), .Q(\mem[27] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i4 (.D(data[3]), .CK(mem_27__7__N_184), .Q(\mem[27] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i5 (.D(data[4]), .CK(mem_27__7__N_184), .Q(\mem[27] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i6 (.D(data[5]), .CK(mem_27__7__N_184), .Q(\mem[27] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i7 (.D(data[6]), .CK(mem_27__7__N_184), .Q(\mem[27] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i8 (.D(data[7]), .CK(mem_27__7__N_184), .Q(\mem[27] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i2 (.D(data[1]), .CK(mem_26__7__N_181), .Q(\mem[26] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i3 (.D(data[2]), .CK(mem_26__7__N_181), .Q(\mem[26] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i4 (.D(data[3]), .CK(mem_26__7__N_181), .Q(\mem[26] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i5 (.D(data[4]), .CK(mem_26__7__N_181), .Q(\mem[26] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i6 (.D(data[5]), .CK(mem_26__7__N_181), .Q(\mem[26] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i7 (.D(data[6]), .CK(mem_26__7__N_181), .Q(\mem[26] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i8 (.D(data[7]), .CK(mem_26__7__N_181), .Q(\mem[26] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i2 (.D(data[1]), .CK(mem_25__7__N_178), .Q(\mem[25] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i3 (.D(data[2]), .CK(mem_25__7__N_178), .Q(\mem[25] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i4 (.D(data[3]), .CK(mem_25__7__N_178), .Q(\mem[25] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i5 (.D(data[4]), .CK(mem_25__7__N_178), .Q(\mem[25] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i6 (.D(data[5]), .CK(mem_25__7__N_178), .Q(\mem[25] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i7 (.D(data[6]), .CK(mem_25__7__N_178), .Q(\mem[25] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i8 (.D(data[7]), .CK(mem_25__7__N_178), .Q(\mem[25] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i2 (.D(data[1]), .CK(mem_24__7__N_175), .Q(\mem[24] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i3 (.D(data[2]), .CK(mem_24__7__N_175), .Q(\mem[24] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i4 (.D(data[3]), .CK(mem_24__7__N_175), .Q(\mem[24] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i5 (.D(data[4]), .CK(mem_24__7__N_175), .Q(\mem[24] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i6 (.D(data[5]), .CK(mem_24__7__N_175), .Q(\mem[24] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i7 (.D(data[6]), .CK(mem_24__7__N_175), .Q(\mem[24] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i8 (.D(data[7]), .CK(mem_24__7__N_175), .Q(\mem[24] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i2 (.D(data[1]), .CK(mem_23__7__N_172), .Q(\mem[23] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i3 (.D(data[2]), .CK(mem_23__7__N_172), .Q(\mem[23] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i4 (.D(data[3]), .CK(mem_23__7__N_172), .Q(\mem[23] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i5 (.D(data[4]), .CK(mem_23__7__N_172), .Q(\mem[23] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i6 (.D(data[5]), .CK(mem_23__7__N_172), .Q(\mem[23] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i7 (.D(data[6]), .CK(mem_23__7__N_172), .Q(\mem[23] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i8 (.D(data[7]), .CK(mem_23__7__N_172), .Q(\mem[23] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i2 (.D(data[1]), .CK(mem_22__7__N_169), .Q(\mem[22] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i3 (.D(data[2]), .CK(mem_22__7__N_169), .Q(\mem[22] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i4 (.D(data[3]), .CK(mem_22__7__N_169), .Q(\mem[22] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i5 (.D(data[4]), .CK(mem_22__7__N_169), .Q(\mem[22] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i6 (.D(data[5]), .CK(mem_22__7__N_169), .Q(\mem[22] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i7 (.D(data[6]), .CK(mem_22__7__N_169), .Q(\mem[22] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i8 (.D(data[7]), .CK(mem_22__7__N_169), .Q(\mem[22] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i2 (.D(data[1]), .CK(mem_21__7__N_166), .Q(\mem[21] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i3 (.D(data[2]), .CK(mem_21__7__N_166), .Q(\mem[21] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i4 (.D(data[3]), .CK(mem_21__7__N_166), .Q(\mem[21] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i5 (.D(data[4]), .CK(mem_21__7__N_166), .Q(\mem[21] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i6 (.D(data[5]), .CK(mem_21__7__N_166), .Q(\mem[21] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i7 (.D(data[6]), .CK(mem_21__7__N_166), .Q(\mem[21] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i8 (.D(data[7]), .CK(mem_21__7__N_166), .Q(\mem[21] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5061_i2 (.D(data[1]), .CK(mem_20__7__N_163), .Q(\mem[20] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5061_i3 (.D(data[2]), .CK(mem_20__7__N_163), .Q(\mem[20] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5061_i4 (.D(data[3]), .CK(mem_20__7__N_163), .Q(\mem[20] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5061_i5 (.D(data[4]), .CK(mem_20__7__N_163), .Q(\mem[20] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5061_i6 (.D(data[5]), .CK(mem_20__7__N_163), .Q(\mem[20] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5061_i7 (.D(data[6]), .CK(mem_20__7__N_163), .Q(\mem[20] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5061_i8 (.D(data[7]), .CK(mem_20__7__N_163), .Q(\mem[20] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i2 (.D(data[1]), .CK(mem_19__7__N_160), .Q(\mem[19] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i3 (.D(data[2]), .CK(mem_19__7__N_160), .Q(\mem[19] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i4 (.D(data[3]), .CK(mem_19__7__N_160), .Q(\mem[19] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i5 (.D(data[4]), .CK(mem_19__7__N_160), .Q(\mem[19] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i6 (.D(data[5]), .CK(mem_19__7__N_160), .Q(\mem[19] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i7 (.D(data[6]), .CK(mem_19__7__N_160), .Q(\mem[19] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i8 (.D(data[7]), .CK(mem_19__7__N_160), .Q(\mem[19] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5055_i2 (.D(data[1]), .CK(mem_18__7__N_157), .Q(\mem[18] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5055_i3 (.D(data[2]), .CK(mem_18__7__N_157), .Q(\mem[18] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5055_i4 (.D(data[3]), .CK(mem_18__7__N_157), .Q(\mem[18] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5055_i5 (.D(data[4]), .CK(mem_18__7__N_157), .Q(\mem[18] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5055_i6 (.D(data[5]), .CK(mem_18__7__N_157), .Q(\mem[18] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5055_i7 (.D(data[6]), .CK(mem_18__7__N_157), .Q(\mem[18] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5055_i8 (.D(data[7]), .CK(mem_18__7__N_157), .Q(\mem[18] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5052_i2 (.D(data[1]), .CK(mem_17__7__N_154), .Q(\mem[17] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5052_i3 (.D(data[2]), .CK(mem_17__7__N_154), .Q(\mem[17] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5052_i4 (.D(data[3]), .CK(mem_17__7__N_154), .Q(\mem[17] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5052_i5 (.D(data[4]), .CK(mem_17__7__N_154), .Q(\mem[17] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5052_i6 (.D(data[5]), .CK(mem_17__7__N_154), .Q(\mem[17] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5052_i7 (.D(data[6]), .CK(mem_17__7__N_154), .Q(\mem[17] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5052_i8 (.D(data[7]), .CK(mem_17__7__N_154), .Q(\mem[17] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i2 (.D(data[1]), .CK(mem_16__7__N_151), .Q(\mem[16] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i3 (.D(data[2]), .CK(mem_16__7__N_151), .Q(\mem[16] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i4 (.D(data[3]), .CK(mem_16__7__N_151), .Q(\mem[16] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i5 (.D(data[4]), .CK(mem_16__7__N_151), .Q(\mem[16] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i6 (.D(data[5]), .CK(mem_16__7__N_151), .Q(\mem[16] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i7 (.D(data[6]), .CK(mem_16__7__N_151), .Q(\mem[16] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i8 (.D(data[7]), .CK(mem_16__7__N_151), .Q(\mem[16] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5046_i2 (.D(data[1]), .CK(mem_15__7__N_148), .Q(\mem[15] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5046_i3 (.D(data[2]), .CK(mem_15__7__N_148), .Q(\mem[15] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5046_i4 (.D(data[3]), .CK(mem_15__7__N_148), .Q(\mem[15] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5046_i5 (.D(data[4]), .CK(mem_15__7__N_148), .Q(\mem[15] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5046_i6 (.D(data[5]), .CK(mem_15__7__N_148), .Q(\mem[15] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5046_i7 (.D(data[6]), .CK(mem_15__7__N_148), .Q(\mem[15] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5046_i8 (.D(data[7]), .CK(mem_15__7__N_148), .Q(\mem[15] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5043_i2 (.D(data[1]), .CK(mem_14__7__N_145), .Q(\mem[14] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5043_i3 (.D(data[2]), .CK(mem_14__7__N_145), .Q(\mem[14] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5043_i4 (.D(data[3]), .CK(mem_14__7__N_145), .Q(\mem[14] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5043_i5 (.D(data[4]), .CK(mem_14__7__N_145), .Q(\mem[14] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5043_i6 (.D(data[5]), .CK(mem_14__7__N_145), .Q(\mem[14] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5043_i7 (.D(data[6]), .CK(mem_14__7__N_145), .Q(\mem[14] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5043_i8 (.D(data[7]), .CK(mem_14__7__N_145), .Q(\mem[14] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5040_i2 (.D(data[1]), .CK(mem_13__7__N_142), .Q(\mem[13] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5040_i3 (.D(data[2]), .CK(mem_13__7__N_142), .Q(\mem[13] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5040_i4 (.D(data[3]), .CK(mem_13__7__N_142), .Q(\mem[13] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5040_i5 (.D(data[4]), .CK(mem_13__7__N_142), .Q(\mem[13] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5040_i6 (.D(data[5]), .CK(mem_13__7__N_142), .Q(\mem[13] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5040_i7 (.D(data[6]), .CK(mem_13__7__N_142), .Q(\mem[13] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5040_i8 (.D(data[7]), .CK(mem_13__7__N_142), .Q(\mem[13] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5037_i2 (.D(data[1]), .CK(mem_12__7__N_139), .Q(\mem[12] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5037_i3 (.D(data[2]), .CK(mem_12__7__N_139), .Q(\mem[12] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5037_i4 (.D(data[3]), .CK(mem_12__7__N_139), .Q(\mem[12] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5037_i5 (.D(data[4]), .CK(mem_12__7__N_139), .Q(\mem[12] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5037_i6 (.D(data[5]), .CK(mem_12__7__N_139), .Q(\mem[12] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5037_i7 (.D(data[6]), .CK(mem_12__7__N_139), .Q(\mem[12] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5037_i8 (.D(data[7]), .CK(mem_12__7__N_139), .Q(\mem[12] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i2 (.D(data[1]), .CK(mem_11__7__N_136), .Q(\mem[11] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i3 (.D(data[2]), .CK(mem_11__7__N_136), .Q(\mem[11] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i4 (.D(data[3]), .CK(mem_11__7__N_136), .Q(\mem[11] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i5 (.D(data[4]), .CK(mem_11__7__N_136), .Q(\mem[11] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i6 (.D(data[5]), .CK(mem_11__7__N_136), .Q(\mem[11] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i7 (.D(data[6]), .CK(mem_11__7__N_136), .Q(\mem[11] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i8 (.D(data[7]), .CK(mem_11__7__N_136), .Q(\mem[11] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5031_i2 (.D(data[1]), .CK(mem_10__7__N_133), .Q(\mem[10] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5031_i3 (.D(data[2]), .CK(mem_10__7__N_133), .Q(\mem[10] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5031_i4 (.D(data[3]), .CK(mem_10__7__N_133), .Q(\mem[10] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5031_i5 (.D(data[4]), .CK(mem_10__7__N_133), .Q(\mem[10] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5031_i6 (.D(data[5]), .CK(mem_10__7__N_133), .Q(\mem[10] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5031_i7 (.D(data[6]), .CK(mem_10__7__N_133), .Q(\mem[10] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5031_i8 (.D(data[7]), .CK(mem_10__7__N_133), .Q(\mem[10] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5028_i2 (.D(data[1]), .CK(mem_9__7__N_130), .Q(\mem[9] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5028_i3 (.D(data[2]), .CK(mem_9__7__N_130), .Q(\mem[9] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5028_i4 (.D(data[3]), .CK(mem_9__7__N_130), .Q(\mem[9] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5028_i5 (.D(data[4]), .CK(mem_9__7__N_130), .Q(\mem[9] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5028_i6 (.D(data[5]), .CK(mem_9__7__N_130), .Q(\mem[9] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5028_i7 (.D(data[6]), .CK(mem_9__7__N_130), .Q(\mem[9] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5028_i8 (.D(data[7]), .CK(mem_9__7__N_130), .Q(\mem[9] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5025_i2 (.D(data[1]), .CK(mem_8__7__N_127), .Q(\mem[8] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5025_i3 (.D(data[2]), .CK(mem_8__7__N_127), .Q(\mem[8] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5025_i4 (.D(data[3]), .CK(mem_8__7__N_127), .Q(\mem[8] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5025_i5 (.D(data[4]), .CK(mem_8__7__N_127), .Q(\mem[8] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5025_i6 (.D(data[5]), .CK(mem_8__7__N_127), .Q(\mem[8] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5025_i7 (.D(data[6]), .CK(mem_8__7__N_127), .Q(\mem[8] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5025_i8 (.D(data[7]), .CK(mem_8__7__N_127), .Q(\mem[8] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5022_i2 (.D(data[1]), .CK(mem_7__7__N_124), .Q(\mem[7] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5022_i3 (.D(data[2]), .CK(mem_7__7__N_124), .Q(\mem[7] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5022_i4 (.D(data[3]), .CK(mem_7__7__N_124), .Q(\mem[7] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5022_i5 (.D(data[4]), .CK(mem_7__7__N_124), .Q(\mem[7] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5022_i6 (.D(data[5]), .CK(mem_7__7__N_124), .Q(\mem[7] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5022_i7 (.D(data[6]), .CK(mem_7__7__N_124), .Q(\mem[7] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5022_i8 (.D(data[7]), .CK(mem_7__7__N_124), .Q(\mem[7] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5019_i2 (.D(data[1]), .CK(mem_6__7__N_121), .Q(\mem[6] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5019_i3 (.D(data[2]), .CK(mem_6__7__N_121), .Q(\mem[6] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5019_i4 (.D(data[3]), .CK(mem_6__7__N_121), .Q(\mem[6] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5019_i5 (.D(data[4]), .CK(mem_6__7__N_121), .Q(\mem[6] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5019_i6 (.D(data[5]), .CK(mem_6__7__N_121), .Q(\mem[6] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5019_i7 (.D(data[6]), .CK(mem_6__7__N_121), .Q(\mem[6] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5019_i8 (.D(data[7]), .CK(mem_6__7__N_121), .Q(\mem[6] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5016_i2 (.D(data[1]), .CK(mem_5__7__N_118), .Q(\mem[5] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5016_i3 (.D(data[2]), .CK(mem_5__7__N_118), .Q(\mem[5] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5016_i4 (.D(data[3]), .CK(mem_5__7__N_118), .Q(\mem[5] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5016_i5 (.D(data[4]), .CK(mem_5__7__N_118), .Q(\mem[5] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5016_i6 (.D(data[5]), .CK(mem_5__7__N_118), .Q(\mem[5] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5016_i7 (.D(data[6]), .CK(mem_5__7__N_118), .Q(\mem[5] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5016_i8 (.D(data[7]), .CK(mem_5__7__N_118), .Q(\mem[5] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i8.GSR = "DISABLED";
    LUT4 i1278_3_lut (.A(\mem[8] [4]), .B(\mem[9] [4]), .C(address[0]), 
         .Z(n1464)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1278_3_lut.init = 16'hcaca;
    LUT4 i1279_3_lut (.A(\mem[10] [4]), .B(\mem[11] [4]), .C(address[0]), 
         .Z(n1465)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1279_3_lut.init = 16'hcaca;
    LUT4 i1280_3_lut (.A(\mem[12] [4]), .B(\mem[13] [4]), .C(address[0]), 
         .Z(n1466)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1280_3_lut.init = 16'hcaca;
    LUT4 i1382_3_lut (.A(\mem[30] [1]), .B(\mem[31] [1]), .C(address[0]), 
         .Z(n1568)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1382_3_lut.init = 16'hcaca;
    LUT4 i1281_3_lut (.A(\mem[14] [4]), .B(\mem[15] [4]), .C(address[0]), 
         .Z(n1467)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1281_3_lut.init = 16'hcaca;
    LUT4 i1282_3_lut (.A(\mem[16] [4]), .B(\mem[17] [4]), .C(address[0]), 
         .Z(n1468)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1282_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_64 (.A(data[7]), .B(akku_o_c_8), .Z(n1895)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_64.init = 16'h8888;
    PFUMX i1512 (.BLUT(n1687), .ALUT(n1688), .C0(address[1]), .Z(n1698));
    LUT4 i893_3_lut_4_lut_4_lut (.A(data[7]), .B(akku_o_c_8), .C(data[5]), 
         .D(data[6]), .Z(\states_2__N_71[2] )) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i893_3_lut_4_lut_4_lut.init = 16'ha8a0;
    LUT4 i1283_3_lut (.A(\mem[18] [4]), .B(\mem[19] [4]), .C(address[0]), 
         .Z(n1469)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1283_3_lut.init = 16'hcaca;
    LUT4 i1284_3_lut (.A(\mem[20] [4]), .B(\mem[21] [4]), .C(address[0]), 
         .Z(n1470)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1284_3_lut.init = 16'hcaca;
    LUT4 i1285_3_lut (.A(\mem[22] [4]), .B(\mem[23] [4]), .C(address[0]), 
         .Z(n1471)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1285_3_lut.init = 16'hcaca;
    LUT4 i1286_3_lut (.A(\mem[24] [4]), .B(\mem[25] [4]), .C(address[0]), 
         .Z(n1472)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1286_3_lut.init = 16'hcaca;
    PFUMX i1513 (.BLUT(n1689), .ALUT(n1690), .C0(address[1]), .Z(n1699));
    LUT4 i1287_3_lut (.A(\mem[26] [4]), .B(\mem[27] [4]), .C(address[0]), 
         .Z(n1473)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1287_3_lut.init = 16'hcaca;
    LUT4 i1381_3_lut (.A(\mem[28] [1]), .B(\mem[29] [1]), .C(address[0]), 
         .Z(n1567)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1381_3_lut.init = 16'hcaca;
    LUT4 i1288_3_lut (.A(\mem[28] [4]), .B(\mem[29] [4]), .C(address[0]), 
         .Z(n1474)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1288_3_lut.init = 16'hcaca;
    PFUMX i1514 (.BLUT(n1691), .ALUT(n1692), .C0(address[1]), .Z(n1700));
    LUT4 i899_4_lut_4_lut (.A(data[7]), .B(akku_o_c_8), .C(data[5]), .D(data[6]), 
         .Z(\states_2__N_71[0] )) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A (D))) */ ;
    defparam i899_4_lut_4_lut.init = 16'h085f;
    LUT4 i1289_3_lut (.A(\mem[30] [4]), .B(\mem[31] [4]), .C(address[0]), 
         .Z(n1475)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1289_3_lut.init = 16'hcaca;
    PFUMX i1352 (.BLUT(n1522), .ALUT(n1523), .C0(address[1]), .Z(n1538));
    LUT4 i1615_3_lut (.A(\mem[32] [7]), .B(\mem[33] [7]), .C(address[0]), 
         .Z(n1801)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1615_3_lut.init = 16'hcaca;
    PFUMX i1353 (.BLUT(n1524), .ALUT(n1525), .C0(address[1]), .Z(n1539));
    LUT4 i1616_3_lut (.A(\mem[34] [7]), .B(\mem[35] [7]), .C(address[0]), 
         .Z(n1802)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1616_3_lut.init = 16'hcaca;
    LUT4 i1617_3_lut (.A(\mem[36] [7]), .B(\mem[37] [7]), .C(address[0]), 
         .Z(n1803)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1617_3_lut.init = 16'hcaca;
    PFUMX i1324 (.BLUT(n1497), .ALUT(n1498), .C0(address[1]), .Z(n1510));
    LUT4 i1618_3_lut (.A(\mem[38] [7]), .B(\mem[39] [7]), .C(address[0]), 
         .Z(n1804)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1618_3_lut.init = 16'hcaca;
    LUT4 i1305_3_lut (.A(\mem[0] [3]), .B(\mem[1] [3]), .C(address[0]), 
         .Z(n1491)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1305_3_lut.init = 16'hcaca;
    PFUMX i1354 (.BLUT(n1526), .ALUT(n1527), .C0(address[1]), .Z(n1540));
    PFUMX i1355 (.BLUT(n1528), .ALUT(n1529), .C0(address[1]), .Z(n1541));
    PFUMX i1356 (.BLUT(n1530), .ALUT(n1531), .C0(address[1]), .Z(n1542));
    PFUMX i1636 (.BLUT(n1811), .ALUT(n1812), .C0(address[1]), .Z(n1822));
    PFUMX i1543 (.BLUT(n1718), .ALUT(n1719), .C0(address[1]), .Z(n1729));
    PFUMX i1357 (.BLUT(n1532), .ALUT(n1533), .C0(address[1]), .Z(n1543));
    PFUMX i1358 (.BLUT(n1534), .ALUT(n1535), .C0(address[1]), .Z(n1544));
    LUT4 i1595_3_lut (.A(\mem[54] [2]), .B(\mem[55] [2]), .C(address[0]), 
         .Z(n1781)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1595_3_lut.init = 16'hcaca;
    PFUMX i1540 (.BLUT(n1712), .ALUT(n1713), .C0(address[1]), .Z(n1726));
    PFUMX i1637 (.BLUT(n1813), .ALUT(n1814), .C0(address[1]), .Z(n1823));
    LUT4 i1594_3_lut (.A(\mem[52] [2]), .B(\mem[53] [2]), .C(address[0]), 
         .Z(n1780)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1594_3_lut.init = 16'hcaca;
    PFUMX i1359 (.BLUT(n1536), .ALUT(n1537), .C0(address[1]), .Z(n1545));
    LUT4 i1159_3_lut (.A(\mem[18] [7]), .B(\mem[19] [7]), .C(address[0]), 
         .Z(n1345)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1159_3_lut.init = 16'hcaca;
    PFUMX i1638 (.BLUT(n1815), .ALUT(n1816), .C0(address[1]), .Z(n1824));
    LUT4 i1397_3_lut (.A(n1581), .B(n1582), .C(address[4]), .Z(n1583)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1397_3_lut.init = 16'hcaca;
    LUT4 i1428_3_lut (.A(n1612), .B(n1613), .C(address[4]), .Z(n1614)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1428_3_lut.init = 16'hcaca;
    LUT4 i1158_3_lut (.A(\mem[16] [7]), .B(\mem[17] [7]), .C(address[0]), 
         .Z(n1344)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1158_3_lut.init = 16'hcaca;
    PFUMX i1600 (.BLUT(n1770), .ALUT(n1771), .C0(address[1]), .Z(n1786));
    LUT4 i1366_3_lut (.A(n1550), .B(n1551), .C(address[4]), .Z(n1552)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1366_3_lut.init = 16'hcaca;
    LUT4 i1459_3_lut (.A(n1643), .B(n1644), .C(address[4]), .Z(n1645)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1459_3_lut.init = 16'hcaca;
    PFUMX i1171 (.BLUT(n1346), .ALUT(n1347), .C0(address[1]), .Z(n1357));
    LUT4 i1335_3_lut (.A(n1519), .B(n1520), .C(address[4]), .Z(n1521)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1335_3_lut.init = 16'hcaca;
    LUT4 i1490_3_lut (.A(n1674), .B(n1675), .C(address[4]), .Z(n1676)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1490_3_lut.init = 16'hcaca;
    LUT4 i1304_3_lut (.A(n1488), .B(n1489), .C(address[4]), .Z(n1490)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1304_3_lut.init = 16'hcaca;
    LUT4 i1521_3_lut (.A(n1705), .B(n1706), .C(address[4]), .Z(n1707)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1521_3_lut.init = 16'hcaca;
    LUT4 i1380_3_lut (.A(\mem[26] [1]), .B(\mem[27] [1]), .C(address[0]), 
         .Z(n1566)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1380_3_lut.init = 16'hcaca;
    LUT4 i1273_3_lut (.A(n1457), .B(n1458), .C(address[4]), .Z(n1459)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1273_3_lut.init = 16'hcaca;
    LUT4 i1552_3_lut (.A(n1736), .B(n1737), .C(address[4]), .Z(n1738)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1552_3_lut.init = 16'hcaca;
    LUT4 i1242_3_lut (.A(n1426), .B(n1427), .C(address[4]), .Z(n1428)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1242_3_lut.init = 16'hcaca;
    LUT4 i1583_3_lut (.A(n1767), .B(n1768), .C(address[4]), .Z(n1769)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1583_3_lut.init = 16'hcaca;
    LUT4 i1211_3_lut (.A(n1395), .B(n1396), .C(address[4]), .Z(n1397)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1211_3_lut.init = 16'hcaca;
    LUT4 i1614_3_lut (.A(n1798), .B(n1799), .C(address[4]), .Z(n1800)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1614_3_lut.init = 16'hcaca;
    LUT4 i1180_3_lut (.A(n1364), .B(n1365), .C(address[4]), .Z(n1366)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1180_3_lut.init = 16'hcaca;
    LUT4 i1645_3_lut (.A(n1829), .B(n1830), .C(address[4]), .Z(n1831)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1645_3_lut.init = 16'hcaca;
    PFUMX i1601 (.BLUT(n1772), .ALUT(n1773), .C0(address[1]), .Z(n1787));
    LUT4 i1398_3_lut (.A(\mem[32] [1]), .B(\mem[33] [1]), .C(address[0]), 
         .Z(n1584)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1398_3_lut.init = 16'hcaca;
    LUT4 i1399_3_lut (.A(\mem[34] [1]), .B(\mem[35] [1]), .C(address[0]), 
         .Z(n1585)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1399_3_lut.init = 16'hcaca;
    LUT4 i1536_3_lut (.A(\mem[60] [5]), .B(\mem[61] [5]), .C(address[0]), 
         .Z(n1722)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1536_3_lut.init = 16'hcaca;
    LUT4 i1537_3_lut (.A(\mem[62] [5]), .B(\mem[63] [5]), .C(address[0]), 
         .Z(n1723)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1537_3_lut.init = 16'hcaca;
    LUT4 i1164_3_lut (.A(\mem[28] [7]), .B(\mem[29] [7]), .C(address[0]), 
         .Z(n1350)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1164_3_lut.init = 16'hcaca;
    LUT4 i1165_3_lut (.A(\mem[30] [7]), .B(\mem[31] [7]), .C(address[0]), 
         .Z(n1351)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1165_3_lut.init = 16'hcaca;
    LUT4 i1400_3_lut (.A(\mem[36] [1]), .B(\mem[37] [1]), .C(address[0]), 
         .Z(n1586)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1400_3_lut.init = 16'hcaca;
    LUT4 i1401_3_lut (.A(\mem[38] [1]), .B(\mem[39] [1]), .C(address[0]), 
         .Z(n1587)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1401_3_lut.init = 16'hcaca;
    LUT4 i1402_3_lut (.A(\mem[40] [1]), .B(\mem[41] [1]), .C(address[0]), 
         .Z(n1588)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1402_3_lut.init = 16'hcaca;
    LUT4 i1403_3_lut (.A(\mem[42] [1]), .B(\mem[43] [1]), .C(address[0]), 
         .Z(n1589)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1403_3_lut.init = 16'hcaca;
    LUT4 i1404_3_lut (.A(\mem[44] [1]), .B(\mem[45] [1]), .C(address[0]), 
         .Z(n1590)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1404_3_lut.init = 16'hcaca;
    LUT4 i1405_3_lut (.A(\mem[46] [1]), .B(\mem[47] [1]), .C(address[0]), 
         .Z(n1591)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1405_3_lut.init = 16'hcaca;
    LUT4 i1406_3_lut (.A(\mem[48] [1]), .B(\mem[49] [1]), .C(address[0]), 
         .Z(n1592)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1406_3_lut.init = 16'hcaca;
    LUT4 i1407_3_lut (.A(\mem[50] [1]), .B(\mem[51] [1]), .C(address[0]), 
         .Z(n1593)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1407_3_lut.init = 16'hcaca;
    LUT4 i1408_3_lut (.A(\mem[52] [1]), .B(\mem[53] [1]), .C(address[0]), 
         .Z(n1594)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1408_3_lut.init = 16'hcaca;
    LUT4 i1409_3_lut (.A(\mem[54] [1]), .B(\mem[55] [1]), .C(address[0]), 
         .Z(n1595)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1409_3_lut.init = 16'hcaca;
    LUT4 i1410_3_lut (.A(\mem[56] [1]), .B(\mem[57] [1]), .C(address[0]), 
         .Z(n1596)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1410_3_lut.init = 16'hcaca;
    LUT4 i1411_3_lut (.A(\mem[58] [1]), .B(\mem[59] [1]), .C(address[0]), 
         .Z(n1597)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1411_3_lut.init = 16'hcaca;
    LUT4 i1412_3_lut (.A(\mem[60] [1]), .B(\mem[61] [1]), .C(address[0]), 
         .Z(n1598)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1412_3_lut.init = 16'hcaca;
    LUT4 i1413_3_lut (.A(\mem[62] [1]), .B(\mem[63] [1]), .C(address[0]), 
         .Z(n1599)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1413_3_lut.init = 16'hcaca;
    LUT4 i1181_3_lut (.A(\mem[0] [2]), .B(\mem[1] [2]), .C(address[0]), 
         .Z(n1367)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1181_3_lut.init = 16'hcaca;
    LUT4 i1182_3_lut (.A(\mem[2] [2]), .B(\mem[3] [2]), .C(address[0]), 
         .Z(n1368)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1182_3_lut.init = 16'hcaca;
    LUT4 i1183_3_lut (.A(\mem[4] [2]), .B(\mem[5] [2]), .C(address[0]), 
         .Z(n1369)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1183_3_lut.init = 16'hcaca;
    LUT4 i1184_3_lut (.A(\mem[6] [2]), .B(\mem[7] [2]), .C(address[0]), 
         .Z(n1370)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1184_3_lut.init = 16'hcaca;
    LUT4 i1185_3_lut (.A(\mem[8] [2]), .B(\mem[9] [2]), .C(address[0]), 
         .Z(n1371)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1185_3_lut.init = 16'hcaca;
    LUT4 i1186_3_lut (.A(\mem[10] [2]), .B(\mem[11] [2]), .C(address[0]), 
         .Z(n1372)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1186_3_lut.init = 16'hcaca;
    LUT4 i1187_3_lut (.A(\mem[12] [2]), .B(\mem[13] [2]), .C(address[0]), 
         .Z(n1373)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1187_3_lut.init = 16'hcaca;
    PFUMX i1602 (.BLUT(n1774), .ALUT(n1775), .C0(address[1]), .Z(n1788));
    LUT4 i1188_3_lut (.A(\mem[14] [2]), .B(\mem[15] [2]), .C(address[0]), 
         .Z(n1374)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1188_3_lut.init = 16'hcaca;
    LUT4 i1189_3_lut (.A(\mem[16] [2]), .B(\mem[17] [2]), .C(address[0]), 
         .Z(n1375)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1189_3_lut.init = 16'hcaca;
    LUT4 i1190_3_lut (.A(\mem[18] [2]), .B(\mem[19] [2]), .C(address[0]), 
         .Z(n1376)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1190_3_lut.init = 16'hcaca;
    LUT4 i1191_3_lut (.A(\mem[20] [2]), .B(\mem[21] [2]), .C(address[0]), 
         .Z(n1377)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1191_3_lut.init = 16'hcaca;
    LUT4 i1192_3_lut (.A(\mem[22] [2]), .B(\mem[23] [2]), .C(address[0]), 
         .Z(n1378)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1192_3_lut.init = 16'hcaca;
    LUT4 i1193_3_lut (.A(\mem[24] [2]), .B(\mem[25] [2]), .C(address[0]), 
         .Z(n1379)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1193_3_lut.init = 16'hcaca;
    LUT4 i1194_3_lut (.A(\mem[26] [2]), .B(\mem[27] [2]), .C(address[0]), 
         .Z(n1380)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1194_3_lut.init = 16'hcaca;
    LUT4 i1195_3_lut (.A(\mem[28] [2]), .B(\mem[29] [2]), .C(address[0]), 
         .Z(n1381)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1195_3_lut.init = 16'hcaca;
    LUT4 i1196_3_lut (.A(\mem[30] [2]), .B(\mem[31] [2]), .C(address[0]), 
         .Z(n1382)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1196_3_lut.init = 16'hcaca;
    LUT4 i1429_3_lut (.A(\mem[32] [0]), .B(\mem[33] [0]), .C(address[0]), 
         .Z(n1615)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1429_3_lut.init = 16'hcaca;
    LUT4 i1430_3_lut (.A(\mem[34] [0]), .B(\mem[35] [0]), .C(address[0]), 
         .Z(n1616)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1430_3_lut.init = 16'hcaca;
    LUT4 i1431_3_lut (.A(\mem[36] [0]), .B(\mem[37] [0]), .C(address[0]), 
         .Z(n1617)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1431_3_lut.init = 16'hcaca;
    LUT4 i1432_3_lut (.A(\mem[38] [0]), .B(\mem[39] [0]), .C(address[0]), 
         .Z(n1618)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1432_3_lut.init = 16'hcaca;
    LUT4 i1433_3_lut (.A(\mem[40] [0]), .B(\mem[41] [0]), .C(address[0]), 
         .Z(n1619)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1433_3_lut.init = 16'hcaca;
    LUT4 i1434_3_lut (.A(\mem[42] [0]), .B(\mem[43] [0]), .C(address[0]), 
         .Z(n1620)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1434_3_lut.init = 16'hcaca;
    LUT4 i1435_3_lut (.A(\mem[44] [0]), .B(\mem[45] [0]), .C(address[0]), 
         .Z(n1621)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1435_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut (.A(address[1]), .B(address[2]), .C(address[0]), .Z(n1302)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i2_3_lut.init = 16'hfbfb;
    LUT4 i1436_3_lut (.A(\mem[46] [0]), .B(\mem[47] [0]), .C(address[0]), 
         .Z(n1622)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1436_3_lut.init = 16'hcaca;
    LUT4 i1437_3_lut (.A(\mem[48] [0]), .B(\mem[49] [0]), .C(address[0]), 
         .Z(n1623)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1437_3_lut.init = 16'hcaca;
    LUT4 i1438_3_lut (.A(\mem[50] [0]), .B(\mem[51] [0]), .C(address[0]), 
         .Z(n1624)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1438_3_lut.init = 16'hcaca;
    LUT4 i1439_3_lut (.A(\mem[52] [0]), .B(\mem[53] [0]), .C(address[0]), 
         .Z(n1625)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1439_3_lut.init = 16'hcaca;
    LUT4 i1440_3_lut (.A(\mem[54] [0]), .B(\mem[55] [0]), .C(address[0]), 
         .Z(n1626)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1440_3_lut.init = 16'hcaca;
    LUT4 i1441_3_lut (.A(\mem[56] [0]), .B(\mem[57] [0]), .C(address[0]), 
         .Z(n1627)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1441_3_lut.init = 16'hcaca;
    LUT4 i1442_3_lut (.A(\mem[58] [0]), .B(\mem[59] [0]), .C(address[0]), 
         .Z(n1628)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1442_3_lut.init = 16'hcaca;
    LUT4 i1443_3_lut (.A(\mem[60] [0]), .B(\mem[61] [0]), .C(address[0]), 
         .Z(n1629)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1443_3_lut.init = 16'hcaca;
    LUT4 i1444_3_lut (.A(\mem[62] [0]), .B(\mem[63] [0]), .C(address[0]), 
         .Z(n1630)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1444_3_lut.init = 16'hcaca;
    LUT4 i1379_3_lut (.A(\mem[24] [1]), .B(\mem[25] [1]), .C(address[0]), 
         .Z(n1565)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1379_3_lut.init = 16'hcaca;
    PFUMX i1603 (.BLUT(n1776), .ALUT(n1777), .C0(address[1]), .Z(n1789));
    LUT4 i1212_3_lut (.A(\mem[0] [6]), .B(\mem[1] [6]), .C(address[0]), 
         .Z(n1398)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1212_3_lut.init = 16'hcaca;
    LUT4 i1213_3_lut (.A(\mem[2] [6]), .B(\mem[3] [6]), .C(address[0]), 
         .Z(n1399)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1213_3_lut.init = 16'hcaca;
    LUT4 i1214_3_lut (.A(\mem[4] [6]), .B(\mem[5] [6]), .C(address[0]), 
         .Z(n1400)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1214_3_lut.init = 16'hcaca;
    LUT4 i1215_3_lut (.A(\mem[6] [6]), .B(\mem[7] [6]), .C(address[0]), 
         .Z(n1401)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1215_3_lut.init = 16'hcaca;
    LUT4 i1216_3_lut (.A(\mem[8] [6]), .B(\mem[9] [6]), .C(address[0]), 
         .Z(n1402)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1216_3_lut.init = 16'hcaca;
    LUT4 i1217_3_lut (.A(\mem[10] [6]), .B(\mem[11] [6]), .C(address[0]), 
         .Z(n1403)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1217_3_lut.init = 16'hcaca;
    LUT4 i1218_3_lut (.A(\mem[12] [6]), .B(\mem[13] [6]), .C(address[0]), 
         .Z(n1404)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1218_3_lut.init = 16'hcaca;
    LUT4 i1219_3_lut (.A(\mem[14] [6]), .B(\mem[15] [6]), .C(address[0]), 
         .Z(n1405)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1219_3_lut.init = 16'hcaca;
    LUT4 i1220_3_lut (.A(\mem[16] [6]), .B(\mem[17] [6]), .C(address[0]), 
         .Z(n1406)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1220_3_lut.init = 16'hcaca;
    LUT4 i1221_3_lut (.A(\mem[18] [6]), .B(\mem[19] [6]), .C(address[0]), 
         .Z(n1407)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1221_3_lut.init = 16'hcaca;
    LUT4 i1222_3_lut (.A(\mem[20] [6]), .B(\mem[21] [6]), .C(address[0]), 
         .Z(n1408)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1222_3_lut.init = 16'hcaca;
    LUT4 i1223_3_lut (.A(\mem[22] [6]), .B(\mem[23] [6]), .C(address[0]), 
         .Z(n1409)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1223_3_lut.init = 16'hcaca;
    LUT4 i1224_3_lut (.A(\mem[24] [6]), .B(\mem[25] [6]), .C(address[0]), 
         .Z(n1410)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1224_3_lut.init = 16'hcaca;
    LUT4 i1225_3_lut (.A(\mem[26] [6]), .B(\mem[27] [6]), .C(address[0]), 
         .Z(n1411)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1225_3_lut.init = 16'hcaca;
    LUT4 i1226_3_lut (.A(\mem[28] [6]), .B(\mem[29] [6]), .C(address[0]), 
         .Z(n1412)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1226_3_lut.init = 16'hcaca;
    LUT4 i1227_3_lut (.A(\mem[30] [6]), .B(\mem[31] [6]), .C(address[0]), 
         .Z(n1413)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1227_3_lut.init = 16'hcaca;
    LUT4 i1553_3_lut (.A(\mem[32] [6]), .B(\mem[33] [6]), .C(address[0]), 
         .Z(n1739)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1553_3_lut.init = 16'hcaca;
    LUT4 i1531_3_lut (.A(\mem[50] [5]), .B(\mem[51] [5]), .C(address[0]), 
         .Z(n1717)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1531_3_lut.init = 16'hcaca;
    PFUMX i1383 (.BLUT(n1553), .ALUT(n1554), .C0(address[1]), .Z(n1569));
    LUT4 i1554_3_lut (.A(\mem[34] [6]), .B(\mem[35] [6]), .C(address[0]), 
         .Z(n1740)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1554_3_lut.init = 16'hcaca;
    LUT4 i1555_3_lut (.A(\mem[36] [6]), .B(\mem[37] [6]), .C(address[0]), 
         .Z(n1741)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1555_3_lut.init = 16'hcaca;
    LUT4 i1556_3_lut (.A(\mem[38] [6]), .B(\mem[39] [6]), .C(address[0]), 
         .Z(n1742)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1556_3_lut.init = 16'hcaca;
    LUT4 i1557_3_lut (.A(\mem[40] [6]), .B(\mem[41] [6]), .C(address[0]), 
         .Z(n1743)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1557_3_lut.init = 16'hcaca;
    LUT4 i1558_3_lut (.A(\mem[42] [6]), .B(\mem[43] [6]), .C(address[0]), 
         .Z(n1744)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1558_3_lut.init = 16'hcaca;
    LUT4 i1243_3_lut (.A(\mem[0] [5]), .B(\mem[1] [5]), .C(address[0]), 
         .Z(n1429)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1243_3_lut.init = 16'hcaca;
    PFUMX i1544 (.BLUT(n1720), .ALUT(n1721), .C0(address[1]), .Z(n1730));
    LUT4 i1244_3_lut (.A(\mem[2] [5]), .B(\mem[3] [5]), .C(address[0]), 
         .Z(n1430)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1244_3_lut.init = 16'hcaca;
    LUT4 i1245_3_lut (.A(\mem[4] [5]), .B(\mem[5] [5]), .C(address[0]), 
         .Z(n1431)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1245_3_lut.init = 16'hcaca;
    LUT4 i1246_3_lut (.A(\mem[6] [5]), .B(\mem[7] [5]), .C(address[0]), 
         .Z(n1432)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1246_3_lut.init = 16'hcaca;
    LUT4 i1559_3_lut (.A(\mem[44] [6]), .B(\mem[45] [6]), .C(address[0]), 
         .Z(n1745)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1559_3_lut.init = 16'hcaca;
    LUT4 i1560_3_lut (.A(\mem[46] [6]), .B(\mem[47] [6]), .C(address[0]), 
         .Z(n1746)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1560_3_lut.init = 16'hcaca;
    LUT4 i1247_3_lut (.A(\mem[8] [5]), .B(\mem[9] [5]), .C(address[0]), 
         .Z(n1433)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1247_3_lut.init = 16'hcaca;
    LUT4 i1248_3_lut (.A(\mem[10] [5]), .B(\mem[11] [5]), .C(address[0]), 
         .Z(n1434)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1248_3_lut.init = 16'hcaca;
    LUT4 i1249_3_lut (.A(\mem[12] [5]), .B(\mem[13] [5]), .C(address[0]), 
         .Z(n1435)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1249_3_lut.init = 16'hcaca;
    LUT4 i1378_3_lut (.A(\mem[22] [1]), .B(\mem[23] [1]), .C(address[0]), 
         .Z(n1564)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1378_3_lut.init = 16'hcaca;
    PFUMX i1541 (.BLUT(n1714), .ALUT(n1715), .C0(address[1]), .Z(n1727));
    LUT4 i1163_3_lut (.A(\mem[26] [7]), .B(\mem[27] [7]), .C(address[0]), 
         .Z(n1349)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1163_3_lut.init = 16'hcaca;
    LUT4 i1529_3_lut (.A(\mem[46] [5]), .B(\mem[47] [5]), .C(address[0]), 
         .Z(n1715)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1529_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut (.A(address[2]), .B(n1904), .C(n1898), .D(n1896), 
         .Z(mem_1__7__N_106)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i1377_3_lut (.A(\mem[20] [1]), .B(\mem[21] [1]), .C(address[0]), 
         .Z(n1563)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1377_3_lut.init = 16'hcaca;
    PFUMX i1384 (.BLUT(n1555), .ALUT(n1556), .C0(address[1]), .Z(n1570));
    LUT4 i1317_3_lut (.A(\mem[24] [3]), .B(\mem[25] [3]), .C(address[0]), 
         .Z(n1503)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1317_3_lut.init = 16'hcaca;
    LUT4 i1598_3_lut (.A(\mem[60] [2]), .B(\mem[61] [2]), .C(address[0]), 
         .Z(n1784)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1598_3_lut.init = 16'hcaca;
    LUT4 i1316_3_lut (.A(\mem[22] [3]), .B(\mem[23] [3]), .C(address[0]), 
         .Z(n1502)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1316_3_lut.init = 16'hcaca;
    LUT4 i1315_3_lut (.A(\mem[20] [3]), .B(\mem[21] [3]), .C(address[0]), 
         .Z(n1501)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1315_3_lut.init = 16'hcaca;
    LUT4 i1376_3_lut (.A(\mem[18] [1]), .B(\mem[19] [1]), .C(address[0]), 
         .Z(n1562)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1376_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_51 (.A(address[2]), .B(n1904), .C(n1906), 
         .D(n1896), .Z(mem_57__7__N_274)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_51.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_52 (.A(address[2]), .B(n1904), .C(n1902), 
         .D(n1896), .Z(mem_49__7__N_250)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_52.init = 16'h0100;
    LUT4 i1_2_lut_3_lut_4_lut_adj_53 (.A(address[2]), .B(n1904), .C(n1901), 
         .D(n1896), .Z(mem_41__7__N_226)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_53.init = 16'h0100;
    LUT4 i1375_3_lut (.A(\mem[16] [1]), .B(\mem[17] [1]), .C(address[0]), 
         .Z(n1561)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1375_3_lut.init = 16'hcaca;
    LUT4 i1374_3_lut (.A(\mem[14] [1]), .B(\mem[15] [1]), .C(address[0]), 
         .Z(n1560)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1374_3_lut.init = 16'hcaca;
    LUT4 i1373_3_lut (.A(\mem[12] [1]), .B(\mem[13] [1]), .C(address[0]), 
         .Z(n1559)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1373_3_lut.init = 16'hcaca;
    LUT4 i1157_3_lut (.A(\mem[14] [7]), .B(\mem[15] [7]), .C(address[0]), 
         .Z(n1343)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1157_3_lut.init = 16'hcaca;
    LUT4 i1156_3_lut (.A(\mem[12] [7]), .B(\mem[13] [7]), .C(address[0]), 
         .Z(n1342)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1156_3_lut.init = 16'hcaca;
    LUT4 i1155_3_lut (.A(\mem[10] [7]), .B(\mem[11] [7]), .C(address[0]), 
         .Z(n1341)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1155_3_lut.init = 16'hcaca;
    PFUMX i1166 (.BLUT(n1336), .ALUT(n1337), .C0(address[1]), .Z(n1352));
    LUT4 i1_2_lut_rep_67_3_lut (.A(address[4]), .B(address[5]), .C(address[3]), 
         .Z(n1898)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_rep_67_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_54 (.A(address[2]), .B(n1904), .C(n1911), 
         .D(n1896), .Z(mem_33__7__N_202)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_54.init = 16'h0100;
    LUT4 i1154_3_lut (.A(\mem[8] [7]), .B(\mem[9] [7]), .C(address[0]), 
         .Z(n1340)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1154_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_55 (.A(address[4]), .B(address[5]), .C(n787), 
         .D(address[3]), .Z(mem_6__7__N_121)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_55.init = 16'h0010;
    LUT4 i1_2_lut_3_lut_4_lut_adj_56 (.A(address[2]), .B(n1904), .C(n1910), 
         .D(n1896), .Z(mem_25__7__N_178)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_56.init = 16'h0100;
    LUT4 i1_2_lut_rep_68_3_lut (.A(address[4]), .B(address[5]), .C(address[3]), 
         .Z(n1899)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_rep_68_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_3_lut_4_lut_adj_57 (.A(address[4]), .B(address[5]), .C(n787), 
         .D(address[3]), .Z(mem_14__7__N_145)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_57.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_58 (.A(address[2]), .B(n1904), .C(n1900), 
         .D(n1896), .Z(mem_17__7__N_154)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_58.init = 16'h0100;
    LUT4 i1_2_lut_3_lut_4_lut_adj_59 (.A(address[2]), .B(n1904), .C(n1899), 
         .D(n1896), .Z(mem_9__7__N_130)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_59.init = 16'h0100;
    LUT4 i2_3_lut_rep_79 (.A(address[3]), .B(address[4]), .C(address[5]), 
         .Z(n1910)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i2_3_lut_rep_79.init = 16'hf7f7;
    LUT4 i1_2_lut_3_lut_4_lut_adj_60 (.A(address[2]), .B(n1904), .C(n1898), 
         .D(n1896), .Z(mem_5__7__N_118)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_60.init = 16'h0200;
    PFUMX i1385 (.BLUT(n1557), .ALUT(n1558), .C0(address[1]), .Z(n1571));
    LUT4 i1_2_lut_4_lut (.A(address[3]), .B(address[4]), .C(address[5]), 
         .D(n787), .Z(mem_30__7__N_193)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_4_lut.init = 16'h0800;
    LUT4 i2_3_lut_rep_80 (.A(address[4]), .B(address[5]), .C(address[3]), 
         .Z(n1911)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i2_3_lut_rep_80.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_4_lut_adj_61 (.A(address[2]), .B(n1904), .C(n1906), 
         .D(n1896), .Z(mem_61__7__N_286)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_61.init = 16'h2000;
    LUT4 i1_2_lut_4_lut_adj_62 (.A(address[4]), .B(address[5]), .C(address[3]), 
         .D(n787), .Z(mem_38__7__N_217)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_4_lut_adj_62.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_63 (.A(address[2]), .B(n1904), .C(n1902), 
         .D(n1896), .Z(mem_53__7__N_262)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_63.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_64 (.A(address[2]), .B(n1904), .C(n1901), 
         .D(n1896), .Z(mem_45__7__N_238)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_64.init = 16'h0200;
    LUT4 i1_2_lut_rep_69_3_lut (.A(address[3]), .B(address[4]), .C(address[5]), 
         .Z(n1900)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_rep_69_3_lut.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_4_lut_adj_65 (.A(address[2]), .B(n1904), .C(n1911), 
         .D(n1896), .Z(mem_37__7__N_214)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_65.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_66 (.A(address[2]), .B(n1904), .C(n1910), 
         .D(n1896), .Z(mem_29__7__N_190)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_66.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_67 (.A(address[2]), .B(n1904), .C(n1900), 
         .D(n1896), .Z(mem_21__7__N_166)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_67.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_68 (.A(address[2]), .B(n1904), .C(n1899), 
         .D(n1896), .Z(mem_13__7__N_142)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_68.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_69 (.A(address[3]), .B(address[4]), .C(n787), 
         .D(address[5]), .Z(mem_22__7__N_169)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_69.init = 16'h0040;
    LUT4 i1_2_lut_rep_71_3_lut (.A(address[3]), .B(address[4]), .C(address[5]), 
         .Z(n1902)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_rep_71_3_lut.init = 16'hbfbf;
    LUT4 i1593_3_lut (.A(\mem[50] [2]), .B(\mem[51] [2]), .C(address[0]), 
         .Z(n1779)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1593_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_70 (.A(address[3]), .B(address[4]), .C(n787), 
         .D(address[5]), .Z(mem_54__7__N_265)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_70.init = 16'h4000;
    PFUMX i1172 (.BLUT(n1348), .ALUT(n1349), .C0(address[1]), .Z(n1358));
    LUT4 i1592_3_lut (.A(\mem[48] [2]), .B(\mem[49] [2]), .C(address[0]), 
         .Z(n1778)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1592_3_lut.init = 16'hcaca;
    PFUMX i1167 (.BLUT(n1338), .ALUT(n1339), .C0(address[1]), .Z(n1353));
    LUT4 i1162_3_lut (.A(\mem[24] [7]), .B(\mem[25] [7]), .C(address[0]), 
         .Z(n1348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1162_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut (.A(address[2]), .B(address[0]), .C(address[1]), 
         .Z(n1327)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut.init = 16'hefef;
    LUT4 i1153_3_lut (.A(\mem[6] [7]), .B(\mem[7] [7]), .C(address[0]), 
         .Z(n1339)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1153_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_71 (.A(address[2]), .B(address[0]), .C(address[1]), 
         .Z(n1328)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_adj_71.init = 16'hfefe;
    LUT4 i1152_3_lut (.A(\mem[4] [7]), .B(\mem[5] [7]), .C(address[0]), 
         .Z(n1338)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1152_3_lut.init = 16'hcaca;
    PFUMX i1604 (.BLUT(n1778), .ALUT(n1779), .C0(address[1]), .Z(n1790));
    LUT4 i1372_3_lut (.A(\mem[10] [1]), .B(\mem[11] [1]), .C(address[0]), 
         .Z(n1558)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1372_3_lut.init = 16'hcaca;
    LUT4 i1497_3_lut (.A(\mem[44] [4]), .B(\mem[45] [4]), .C(address[0]), 
         .Z(n1683)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1497_3_lut.init = 16'hcaca;
    PFUMX i1168 (.BLUT(n1340), .ALUT(n1341), .C0(address[1]), .Z(n1354));
    LUT4 i1371_3_lut (.A(\mem[8] [1]), .B(\mem[9] [1]), .C(address[0]), 
         .Z(n1557)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1371_3_lut.init = 16'hcaca;
    LUT4 i1624_3_lut (.A(\mem[50] [7]), .B(\mem[51] [7]), .C(address[0]), 
         .Z(n1810)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1624_3_lut.init = 16'hcaca;
    PFUMX i1169 (.BLUT(n1342), .ALUT(n1343), .C0(address[1]), .Z(n1355));
    PFUMX i1386 (.BLUT(n1559), .ALUT(n1560), .C0(address[1]), .Z(n1572));
    LUT4 Select_406_i3_4_lut (.A(data_7__N_84[1]), .B(akku_o_c_1), .C(data_7__N_97), 
         .D(n1905), .Z(data[1])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_406_i3_4_lut.init = 16'ha0ec;
    PFUMX i1387 (.BLUT(n1561), .ALUT(n1562), .C0(address[1]), .Z(n1573));
    LUT4 i1151_3_lut (.A(\mem[2] [7]), .B(\mem[3] [7]), .C(address[0]), 
         .Z(n1337)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1151_3_lut.init = 16'hcaca;
    LUT4 i1150_3_lut (.A(\mem[0] [7]), .B(\mem[1] [7]), .C(address[0]), 
         .Z(n1336)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1150_3_lut.init = 16'hcaca;
    PFUMX i1388 (.BLUT(n1563), .ALUT(n1564), .C0(address[1]), .Z(n1574));
    LUT4 Select_405_i3_4_lut (.A(data_7__N_84[2]), .B(akku_o_c_2), .C(data_7__N_97), 
         .D(n1905), .Z(data[2])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_405_i3_4_lut.init = 16'ha0ec;
    LUT4 Select_404_i3_4_lut (.A(data_7__N_84[3]), .B(akku_o_c_3), .C(data_7__N_97), 
         .D(n1905), .Z(data[3])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_404_i3_4_lut.init = 16'ha0ec;
    LUT4 Select_403_i3_4_lut (.A(data_7__N_84[4]), .B(akku_o_c_4), .C(data_7__N_97), 
         .D(n1905), .Z(data[4])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_403_i3_4_lut.init = 16'ha0ec;
    LUT4 Select_402_i3_4_lut (.A(data_7__N_84[5]), .B(akku_o_c_5), .C(data_7__N_97), 
         .D(n1905), .Z(data[5])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_402_i3_4_lut.init = 16'ha0ec;
    LUT4 Select_401_i3_4_lut (.A(data_7__N_84[6]), .B(akku_o_c_6), .C(data_7__N_97), 
         .D(n1905), .Z(data[6])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_401_i3_4_lut.init = 16'ha0ec;
    LUT4 Select_400_i3_4_lut (.A(data_7__N_84[7]), .B(akku_o_c_7), .C(data_7__N_97), 
         .D(n1905), .Z(data[7])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam Select_400_i3_4_lut.init = 16'ha0ec;
    LUT4 i1370_3_lut (.A(\mem[6] [1]), .B(\mem[7] [1]), .C(address[0]), 
         .Z(n1556)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1370_3_lut.init = 16'hcaca;
    LUT4 i1535_3_lut (.A(\mem[58] [5]), .B(\mem[59] [5]), .C(address[0]), 
         .Z(n1721)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1535_3_lut.init = 16'hcaca;
    LUT4 i1528_3_lut (.A(\mem[44] [5]), .B(\mem[45] [5]), .C(address[0]), 
         .Z(n1714)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1528_3_lut.init = 16'hcaca;
    LUT4 i1369_3_lut (.A(\mem[4] [1]), .B(\mem[5] [1]), .C(address[0]), 
         .Z(n1555)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1369_3_lut.init = 16'hcaca;
    LUT4 i1534_3_lut (.A(\mem[56] [5]), .B(\mem[57] [5]), .C(address[0]), 
         .Z(n1720)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1534_3_lut.init = 16'hcaca;
    LUT4 i1368_3_lut (.A(\mem[2] [1]), .B(\mem[3] [1]), .C(address[0]), 
         .Z(n1554)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1368_3_lut.init = 16'hcaca;
    LUT4 i1367_3_lut (.A(\mem[0] [1]), .B(\mem[1] [1]), .C(address[0]), 
         .Z(n1553)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1367_3_lut.init = 16'hcaca;
    LUT4 i1591_3_lut (.A(\mem[46] [2]), .B(\mem[47] [2]), .C(address[0]), 
         .Z(n1777)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1591_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_70_3_lut (.A(address[5]), .B(address[3]), .C(address[4]), 
         .Z(n1901)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_rep_70_3_lut.init = 16'hf7f7;
    LUT4 i1590_3_lut (.A(\mem[44] [2]), .B(\mem[45] [2]), .C(address[0]), 
         .Z(n1776)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1590_3_lut.init = 16'hcaca;
    LUT4 i1589_3_lut (.A(\mem[42] [2]), .B(\mem[43] [2]), .C(address[0]), 
         .Z(n1775)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1589_3_lut.init = 16'hcaca;
    LUT4 i1588_3_lut (.A(\mem[40] [2]), .B(\mem[41] [2]), .C(address[0]), 
         .Z(n1774)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1588_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_72 (.A(address[5]), .B(address[3]), .C(n787), 
         .D(address[4]), .Z(mem_46__7__N_241)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_72.init = 16'h0080;
    LUT4 i1161_3_lut (.A(\mem[22] [7]), .B(\mem[23] [7]), .C(address[0]), 
         .Z(n1347)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1161_3_lut.init = 16'hcaca;
    LUT4 i1527_3_lut (.A(\mem[42] [5]), .B(\mem[43] [5]), .C(address[0]), 
         .Z(n1713)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1527_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_75_3_lut (.A(address[5]), .B(address[3]), .C(address[4]), 
         .Z(n1906)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_75_3_lut.init = 16'h8080;
    LUT4 i1587_3_lut (.A(\mem[38] [2]), .B(\mem[39] [2]), .C(address[0]), 
         .Z(n1773)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1587_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_73 (.A(address[5]), .B(address[3]), .C(n787), 
         .D(address[4]), .Z(mem_62__7__N_289)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_73.init = 16'h8000;
    LUT4 i1586_3_lut (.A(\mem[36] [2]), .B(\mem[37] [2]), .C(address[0]), 
         .Z(n1772)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1586_3_lut.init = 16'hcaca;
    LUT4 i400_1_lut_rep_85 (.A(address[0]), .Z(n1916)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i400_1_lut_rep_85.init = 16'h5555;
    LUT4 i3_4_lut_4_lut (.A(address[0]), .B(address[1]), .C(address[2]), 
         .D(n1896), .Z(n787)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i3_4_lut_4_lut.init = 16'h4000;
    LUT4 i1160_3_lut (.A(\mem[20] [7]), .B(\mem[21] [7]), .C(address[0]), 
         .Z(n1346)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1160_3_lut.init = 16'hcaca;
    LUT4 i1585_3_lut (.A(\mem[34] [2]), .B(\mem[35] [2]), .C(address[0]), 
         .Z(n1771)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1585_3_lut.init = 16'hcaca;
    LUT4 i1584_3_lut (.A(\mem[32] [2]), .B(\mem[33] [2]), .C(address[0]), 
         .Z(n1770)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1584_3_lut.init = 16'hcaca;
    PFUMX i1389 (.BLUT(n1565), .ALUT(n1566), .C0(address[1]), .Z(n1575));
    LUT4 i1630_3_lut (.A(\mem[62] [7]), .B(\mem[63] [7]), .C(address[0]), 
         .Z(n1816)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1630_3_lut.init = 16'hcaca;
    LUT4 i1629_3_lut (.A(\mem[60] [7]), .B(\mem[61] [7]), .C(address[0]), 
         .Z(n1815)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1629_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_73_2_lut (.A(address[0]), .B(address[1]), .Z(n1904)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_rep_73_2_lut.init = 16'hdddd;
    LUT4 i1351_3_lut (.A(\mem[30] [0]), .B(\mem[31] [0]), .C(address[0]), 
         .Z(n1537)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1351_3_lut.init = 16'hcaca;
    LUT4 i1350_3_lut (.A(\mem[28] [0]), .B(\mem[29] [0]), .C(address[0]), 
         .Z(n1536)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1350_3_lut.init = 16'hcaca;
    LUT4 i1533_3_lut (.A(\mem[54] [5]), .B(\mem[55] [5]), .C(address[0]), 
         .Z(n1719)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1533_3_lut.init = 16'hcaca;
    LUT4 i1526_3_lut (.A(\mem[40] [5]), .B(\mem[41] [5]), .C(address[0]), 
         .Z(n1712)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1526_3_lut.init = 16'hcaca;
    LUT4 i1628_3_lut (.A(\mem[58] [7]), .B(\mem[59] [7]), .C(address[0]), 
         .Z(n1814)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1628_3_lut.init = 16'hcaca;
    LUT4 i1627_3_lut (.A(\mem[56] [7]), .B(\mem[57] [7]), .C(address[0]), 
         .Z(n1813)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1627_3_lut.init = 16'hcaca;
    LUT4 i1532_3_lut (.A(\mem[52] [5]), .B(\mem[53] [5]), .C(address[0]), 
         .Z(n1718)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1532_3_lut.init = 16'hcaca;
    LUT4 i1349_3_lut (.A(\mem[26] [0]), .B(\mem[27] [0]), .C(address[0]), 
         .Z(n1535)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1349_3_lut.init = 16'hcaca;
    LUT4 i1525_3_lut (.A(\mem[38] [5]), .B(\mem[39] [5]), .C(address[0]), 
         .Z(n1711)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1525_3_lut.init = 16'hcaca;
    LUT4 i1348_3_lut (.A(\mem[24] [0]), .B(\mem[25] [0]), .C(address[0]), 
         .Z(n1534)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1348_3_lut.init = 16'hcaca;
    LUT4 i1347_3_lut (.A(\mem[22] [0]), .B(\mem[23] [0]), .C(address[0]), 
         .Z(n1533)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1347_3_lut.init = 16'hcaca;
    LUT4 i1346_3_lut (.A(\mem[20] [0]), .B(\mem[21] [0]), .C(address[0]), 
         .Z(n1532)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1346_3_lut.init = 16'hcaca;
    LUT4 i1626_3_lut (.A(\mem[54] [7]), .B(\mem[55] [7]), .C(address[0]), 
         .Z(n1812)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1626_3_lut.init = 16'hcaca;
    LUT4 i1625_3_lut (.A(\mem[52] [7]), .B(\mem[53] [7]), .C(address[0]), 
         .Z(n1811)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1625_3_lut.init = 16'hcaca;
    PFUMX i1170 (.BLUT(n1344), .ALUT(n1345), .C0(address[1]), .Z(n1356));
    PFUMX i1542 (.BLUT(n1716), .ALUT(n1717), .C0(address[1]), .Z(n1728));
    LUT4 i1345_3_lut (.A(\mem[18] [0]), .B(\mem[19] [0]), .C(address[0]), 
         .Z(n1531)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1345_3_lut.init = 16'hcaca;
    LUT4 i1344_3_lut (.A(\mem[16] [0]), .B(\mem[17] [0]), .C(address[0]), 
         .Z(n1530)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1344_3_lut.init = 16'hcaca;
    LUT4 i1343_3_lut (.A(\mem[14] [0]), .B(\mem[15] [0]), .C(address[0]), 
         .Z(n1529)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1343_3_lut.init = 16'hcaca;
    LUT4 i1342_3_lut (.A(\mem[12] [0]), .B(\mem[13] [0]), .C(address[0]), 
         .Z(n1528)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1342_3_lut.init = 16'hcaca;
    LUT4 i1341_3_lut (.A(\mem[10] [0]), .B(\mem[11] [0]), .C(address[0]), 
         .Z(n1527)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1341_3_lut.init = 16'hcaca;
    LUT4 i1340_3_lut (.A(\mem[8] [0]), .B(\mem[9] [0]), .C(address[0]), 
         .Z(n1526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1340_3_lut.init = 16'hcaca;
    LUT4 i1339_3_lut (.A(\mem[6] [0]), .B(\mem[7] [0]), .C(address[0]), 
         .Z(n1525)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1339_3_lut.init = 16'hcaca;
    LUT4 i1338_3_lut (.A(\mem[4] [0]), .B(\mem[5] [0]), .C(address[0]), 
         .Z(n1524)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1338_3_lut.init = 16'hcaca;
    LUT4 i1337_3_lut (.A(\mem[2] [0]), .B(\mem[3] [0]), .C(address[0]), 
         .Z(n1523)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1337_3_lut.init = 16'hcaca;
    LUT4 i1336_3_lut (.A(\mem[0] [0]), .B(\mem[1] [0]), .C(address[0]), 
         .Z(n1522)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1336_3_lut.init = 16'hcaca;
    LUT4 i1506_3_lut (.A(\mem[62] [4]), .B(\mem[63] [4]), .C(address[0]), 
         .Z(n1692)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1506_3_lut.init = 16'hcaca;
    LUT4 i1505_3_lut (.A(\mem[60] [4]), .B(\mem[61] [4]), .C(address[0]), 
         .Z(n1691)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1505_3_lut.init = 16'hcaca;
    PFUMX i1605 (.BLUT(n1780), .ALUT(n1781), .C0(address[1]), .Z(n1791));
    LUT4 i1311_3_lut (.A(\mem[12] [3]), .B(\mem[13] [3]), .C(address[0]), 
         .Z(n1497)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1311_3_lut.init = 16'hcaca;
    LUT4 i1498_3_lut (.A(\mem[46] [4]), .B(\mem[47] [4]), .C(address[0]), 
         .Z(n1684)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1498_3_lut.init = 16'hcaca;
    LUT4 i1499_3_lut (.A(\mem[48] [4]), .B(\mem[49] [4]), .C(address[0]), 
         .Z(n1685)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1499_3_lut.init = 16'hcaca;
    LUT4 i1500_3_lut (.A(\mem[50] [4]), .B(\mem[51] [4]), .C(address[0]), 
         .Z(n1686)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1500_3_lut.init = 16'hcaca;
    PFUMX i1390 (.BLUT(n1567), .ALUT(n1568), .C0(address[1]), .Z(n1576));
    LUT4 i1504_3_lut (.A(\mem[58] [4]), .B(\mem[59] [4]), .C(address[0]), 
         .Z(n1690)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1504_3_lut.init = 16'hcaca;
    LUT4 i1503_3_lut (.A(\mem[56] [4]), .B(\mem[57] [4]), .C(address[0]), 
         .Z(n1689)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1503_3_lut.init = 16'hcaca;
    LUT4 i1530_3_lut (.A(\mem[48] [5]), .B(\mem[49] [5]), .C(address[0]), 
         .Z(n1716)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1530_3_lut.init = 16'hcaca;
    LUT4 i1623_3_lut (.A(\mem[48] [7]), .B(\mem[49] [7]), .C(address[0]), 
         .Z(n1809)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1623_3_lut.init = 16'hcaca;
    LUT4 i1599_3_lut (.A(\mem[62] [2]), .B(\mem[63] [2]), .C(address[0]), 
         .Z(n1785)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1599_3_lut.init = 16'hcaca;
    LUT4 i1501_3_lut (.A(\mem[52] [4]), .B(\mem[53] [4]), .C(address[0]), 
         .Z(n1687)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1501_3_lut.init = 16'hcaca;
    LUT4 i1622_3_lut (.A(\mem[46] [7]), .B(\mem[47] [7]), .C(address[0]), 
         .Z(n1808)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1622_3_lut.init = 16'hcaca;
    LUT4 i1621_3_lut (.A(\mem[44] [7]), .B(\mem[45] [7]), .C(address[0]), 
         .Z(n1807)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1621_3_lut.init = 16'hcaca;
    LUT4 i1496_3_lut (.A(\mem[42] [4]), .B(\mem[43] [4]), .C(address[0]), 
         .Z(n1682)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1496_3_lut.init = 16'hcaca;
    LUT4 i1495_3_lut (.A(\mem[40] [4]), .B(\mem[41] [4]), .C(address[0]), 
         .Z(n1681)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1495_3_lut.init = 16'hcaca;
    LUT4 i1494_3_lut (.A(\mem[38] [4]), .B(\mem[39] [4]), .C(address[0]), 
         .Z(n1680)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1494_3_lut.init = 16'hcaca;
    LUT4 i1493_3_lut (.A(\mem[36] [4]), .B(\mem[37] [4]), .C(address[0]), 
         .Z(n1679)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1493_3_lut.init = 16'hcaca;
    LUT4 i1492_3_lut (.A(\mem[34] [4]), .B(\mem[35] [4]), .C(address[0]), 
         .Z(n1678)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1492_3_lut.init = 16'hcaca;
    LUT4 i1491_3_lut (.A(\mem[32] [4]), .B(\mem[33] [4]), .C(address[0]), 
         .Z(n1677)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1491_3_lut.init = 16'hcaca;
    LUT4 i1620_3_lut (.A(\mem[42] [7]), .B(\mem[43] [7]), .C(address[0]), 
         .Z(n1806)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1620_3_lut.init = 16'hcaca;
    LUT4 i1619_3_lut (.A(\mem[40] [7]), .B(\mem[41] [7]), .C(address[0]), 
         .Z(n1805)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1619_3_lut.init = 16'hcaca;
    LUT4 i1320_3_lut (.A(\mem[30] [3]), .B(\mem[31] [3]), .C(address[0]), 
         .Z(n1506)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1320_3_lut.init = 16'hcaca;
    LUT4 i1319_3_lut (.A(\mem[28] [3]), .B(\mem[29] [3]), .C(address[0]), 
         .Z(n1505)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1319_3_lut.init = 16'hcaca;
    LUT4 i1318_3_lut (.A(\mem[26] [3]), .B(\mem[27] [3]), .C(address[0]), 
         .Z(n1504)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1318_3_lut.init = 16'hcaca;
    LUT4 i1314_3_lut (.A(\mem[18] [3]), .B(\mem[19] [3]), .C(address[0]), 
         .Z(n1500)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1314_3_lut.init = 16'hcaca;
    PFUMX i1606 (.BLUT(n1782), .ALUT(n1783), .C0(address[1]), .Z(n1792));
    LUT4 i1312_3_lut (.A(\mem[14] [3]), .B(\mem[15] [3]), .C(address[0]), 
         .Z(n1498)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1312_3_lut.init = 16'hcaca;
    LUT4 i1502_3_lut (.A(\mem[54] [4]), .B(\mem[55] [4]), .C(address[0]), 
         .Z(n1688)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i1502_3_lut.init = 16'hcaca;
    PFUMX i1538 (.BLUT(n1708), .ALUT(n1709), .C0(address[1]), .Z(n1724));
    PFUMX i1539 (.BLUT(n1710), .ALUT(n1711), .C0(address[1]), .Z(n1725));
    PFUMX i1325 (.BLUT(n1499), .ALUT(n1500), .C0(address[1]), .Z(n1511));
    PFUMX i1323 (.BLUT(n1495), .ALUT(n1496), .C0(address[1]), .Z(n1509));
    PFUMX i1322 (.BLUT(n1493), .ALUT(n1494), .C0(address[1]), .Z(n1508));
    PFUMX i1321 (.BLUT(n1491), .ALUT(n1492), .C0(address[1]), .Z(n1507));
    PFUMX i1632 (.BLUT(n1803), .ALUT(n1804), .C0(address[1]), .Z(n1818));
    PFUMX i1631 (.BLUT(n1801), .ALUT(n1802), .C0(address[1]), .Z(n1817));
    PFUMX i1297 (.BLUT(n1474), .ALUT(n1475), .C0(address[1]), .Z(n1483));
    PFUMX i1296 (.BLUT(n1472), .ALUT(n1473), .C0(address[1]), .Z(n1482));
    PFUMX i1295 (.BLUT(n1470), .ALUT(n1471), .C0(address[1]), .Z(n1481));
    PFUMX i1294 (.BLUT(n1468), .ALUT(n1469), .C0(address[1]), .Z(n1480));
    PFUMX i1293 (.BLUT(n1466), .ALUT(n1467), .C0(address[1]), .Z(n1479));
    PFUMX i1292 (.BLUT(n1464), .ALUT(n1465), .C0(address[1]), .Z(n1478));
    PFUMX i1291 (.BLUT(n1462), .ALUT(n1463), .C0(address[1]), .Z(n1477));
    PFUMX i1483 (.BLUT(n1660), .ALUT(n1661), .C0(address[1]), .Z(n1669));
    PFUMX i1290 (.BLUT(n1460), .ALUT(n1461), .C0(address[1]), .Z(n1476));
    PFUMX i1482 (.BLUT(n1658), .ALUT(n1659), .C0(address[1]), .Z(n1668));
    PFUMX i1481 (.BLUT(n1656), .ALUT(n1657), .C0(address[1]), .Z(n1667));
    PFUMX i1480 (.BLUT(n1654), .ALUT(n1655), .C0(address[1]), .Z(n1666));
    PFUMX i1479 (.BLUT(n1652), .ALUT(n1653), .C0(address[1]), .Z(n1665));
    PFUMX i1478 (.BLUT(n1650), .ALUT(n1651), .C0(address[1]), .Z(n1664));
    PFUMX i1477 (.BLUT(n1648), .ALUT(n1649), .C0(address[1]), .Z(n1663));
    PFUMX i1576 (.BLUT(n1753), .ALUT(n1754), .C0(address[1]), .Z(n1762));
    PFUMX i1575 (.BLUT(n1751), .ALUT(n1752), .C0(address[1]), .Z(n1761));
    PFUMX i1476 (.BLUT(n1646), .ALUT(n1647), .C0(address[1]), .Z(n1662));
    PFUMX i1574 (.BLUT(n1749), .ALUT(n1750), .C0(address[1]), .Z(n1760));
    PFUMX i1266 (.BLUT(n1443), .ALUT(n1444), .C0(address[1]), .Z(n1452));
    PFUMX i1265 (.BLUT(n1441), .ALUT(n1442), .C0(address[1]), .Z(n1451));
    PFUMX i1573 (.BLUT(n1747), .ALUT(n1748), .C0(address[1]), .Z(n1759));
    PFUMX i1264 (.BLUT(n1439), .ALUT(n1440), .C0(address[1]), .Z(n1450));
    PFUMX i1263 (.BLUT(n1437), .ALUT(n1438), .C0(address[1]), .Z(n1449));
    PFUMX i1262 (.BLUT(n1435), .ALUT(n1436), .C0(address[1]), .Z(n1448));
    PFUMX i1261 (.BLUT(n1433), .ALUT(n1434), .C0(address[1]), .Z(n1447));
    PFUMX i1572 (.BLUT(n1745), .ALUT(n1746), .C0(address[1]), .Z(n1758));
    PFUMX i1260 (.BLUT(n1431), .ALUT(n1432), .C0(address[1]), .Z(n1446));
    PFUMX i1259 (.BLUT(n1429), .ALUT(n1430), .C0(address[1]), .Z(n1445));
    PFUMX i1571 (.BLUT(n1743), .ALUT(n1744), .C0(address[1]), .Z(n1757));
    PFUMX i1570 (.BLUT(n1741), .ALUT(n1742), .C0(address[1]), .Z(n1756));
    PFUMX i1569 (.BLUT(n1739), .ALUT(n1740), .C0(address[1]), .Z(n1755));
    PFUMX i1235 (.BLUT(n1412), .ALUT(n1413), .C0(address[1]), .Z(n1421));
    PFUMX i1234 (.BLUT(n1410), .ALUT(n1411), .C0(address[1]), .Z(n1420));
    PFUMX i1233 (.BLUT(n1408), .ALUT(n1409), .C0(address[1]), .Z(n1419));
    PFUMX i1232 (.BLUT(n1406), .ALUT(n1407), .C0(address[1]), .Z(n1418));
    PFUMX i1231 (.BLUT(n1404), .ALUT(n1405), .C0(address[1]), .Z(n1417));
    PFUMX i1230 (.BLUT(n1402), .ALUT(n1403), .C0(address[1]), .Z(n1416));
    PFUMX i1229 (.BLUT(n1400), .ALUT(n1401), .C0(address[1]), .Z(n1415));
    PFUMX i1228 (.BLUT(n1398), .ALUT(n1399), .C0(address[1]), .Z(n1414));
    PFUMX i1452 (.BLUT(n1629), .ALUT(n1630), .C0(address[1]), .Z(n1638));
    PFUMX i1451 (.BLUT(n1627), .ALUT(n1628), .C0(address[1]), .Z(n1637));
    PFUMX i1450 (.BLUT(n1625), .ALUT(n1626), .C0(address[1]), .Z(n1636));
    PFUMX i1449 (.BLUT(n1623), .ALUT(n1624), .C0(address[1]), .Z(n1635));
    PFUMX i1448 (.BLUT(n1621), .ALUT(n1622), .C0(address[1]), .Z(n1634));
    PFUMX i1447 (.BLUT(n1619), .ALUT(n1620), .C0(address[1]), .Z(n1633));
    PFUMX i1446 (.BLUT(n1617), .ALUT(n1618), .C0(address[1]), .Z(n1632));
    PFUMX i1445 (.BLUT(n1615), .ALUT(n1616), .C0(address[1]), .Z(n1631));
    PFUMX i1204 (.BLUT(n1381), .ALUT(n1382), .C0(address[1]), .Z(n1390));
    PFUMX i1203 (.BLUT(n1379), .ALUT(n1380), .C0(address[1]), .Z(n1389));
    PFUMX i1202 (.BLUT(n1377), .ALUT(n1378), .C0(address[1]), .Z(n1388));
    PFUMX i1201 (.BLUT(n1375), .ALUT(n1376), .C0(address[1]), .Z(n1387));
    PFUMX i1200 (.BLUT(n1373), .ALUT(n1374), .C0(address[1]), .Z(n1386));
    PFUMX i1199 (.BLUT(n1371), .ALUT(n1372), .C0(address[1]), .Z(n1385));
    PFUMX i1198 (.BLUT(n1369), .ALUT(n1370), .C0(address[1]), .Z(n1384));
    PFUMX i1197 (.BLUT(n1367), .ALUT(n1368), .C0(address[1]), .Z(n1383));
    PFUMX i1421 (.BLUT(n1598), .ALUT(n1599), .C0(address[1]), .Z(n1607));
    PFUMX i1420 (.BLUT(n1596), .ALUT(n1597), .C0(address[1]), .Z(n1606));
    PFUMX i1419 (.BLUT(n1594), .ALUT(n1595), .C0(address[1]), .Z(n1605));
    PFUMX i1418 (.BLUT(n1592), .ALUT(n1593), .C0(address[1]), .Z(n1604));
    PFUMX i1417 (.BLUT(n1590), .ALUT(n1591), .C0(address[1]), .Z(n1603));
    PFUMX i1416 (.BLUT(n1588), .ALUT(n1589), .C0(address[1]), .Z(n1602));
    PFUMX i1415 (.BLUT(n1586), .ALUT(n1587), .C0(address[1]), .Z(n1601));
    PFUMX i1173 (.BLUT(n1350), .ALUT(n1351), .C0(address[1]), .Z(n1359));
    PFUMX i1545 (.BLUT(n1722), .ALUT(n1723), .C0(address[1]), .Z(n1731));
    PFUMX i1414 (.BLUT(n1584), .ALUT(n1585), .C0(address[1]), .Z(n1600));
    L6MUX21 i1610 (.D0(n1790), .D1(n1791), .SD(address[2]), .Z(n1796));
    L6MUX21 i1609 (.D0(n1788), .D1(n1789), .SD(address[2]), .Z(n1795));
    L6MUX21 i1642 (.D0(n1823), .D1(n1824), .SD(address[2]), .Z(n1828));
    L6MUX21 i1608 (.D0(n1786), .D1(n1787), .SD(address[2]), .Z(n1794));
    L6MUX21 i1394 (.D0(n1575), .D1(n1576), .SD(address[2]), .Z(n1580));
    L6MUX21 i1393 (.D0(n1573), .D1(n1574), .SD(address[2]), .Z(n1579));
    L6MUX21 i1392 (.D0(n1571), .D1(n1572), .SD(address[2]), .Z(n1578));
    L6MUX21 i1391 (.D0(n1569), .D1(n1570), .SD(address[2]), .Z(n1577));
    L6MUX21 i1641 (.D0(n1821), .D1(n1822), .SD(address[2]), .Z(n1827));
    L6MUX21 i1640 (.D0(n1819), .D1(n1820), .SD(address[2]), .Z(n1826));
    L6MUX21 i1639 (.D0(n1817), .D1(n1818), .SD(address[2]), .Z(n1825));
    L6MUX21 i1363 (.D0(n1544), .D1(n1545), .SD(address[2]), .Z(n1549));
    L6MUX21 i1362 (.D0(n1542), .D1(n1543), .SD(address[2]), .Z(n1548));
    L6MUX21 i1361 (.D0(n1540), .D1(n1541), .SD(address[2]), .Z(n1547));
    L6MUX21 i1360 (.D0(n1538), .D1(n1539), .SD(address[2]), .Z(n1546));
    L6MUX21 i1518 (.D0(n1699), .D1(n1700), .SD(address[2]), .Z(n1704));
    L6MUX21 i1517 (.D0(n1697), .D1(n1698), .SD(address[2]), .Z(n1703));
    L6MUX21 i1516 (.D0(n1695), .D1(n1696), .SD(address[2]), .Z(n1702));
    L6MUX21 i1515 (.D0(n1693), .D1(n1694), .SD(address[2]), .Z(n1701));
    L6MUX21 i1332 (.D0(n1513), .D1(n1514), .SD(address[2]), .Z(n1518));
    L6MUX21 i1331 (.D0(n1511), .D1(n1512), .SD(address[2]), .Z(n1517));
    L6MUX21 i1330 (.D0(n1509), .D1(n1510), .SD(address[2]), .Z(n1516));
    L6MUX21 i1329 (.D0(n1507), .D1(n1508), .SD(address[2]), .Z(n1515));
    L6MUX21 i1301 (.D0(n1482), .D1(n1483), .SD(address[2]), .Z(n1487));
    L6MUX21 i1300 (.D0(n1480), .D1(n1481), .SD(address[2]), .Z(n1486));
    L6MUX21 i1299 (.D0(n1478), .D1(n1479), .SD(address[2]), .Z(n1485));
    L6MUX21 i1298 (.D0(n1476), .D1(n1477), .SD(address[2]), .Z(n1484));
    L6MUX21 i1487 (.D0(n1668), .D1(n1669), .SD(address[2]), .Z(n1673));
    L6MUX21 i1486 (.D0(n1666), .D1(n1667), .SD(address[2]), .Z(n1672));
    L6MUX21 i1485 (.D0(n1664), .D1(n1665), .SD(address[2]), .Z(n1671));
    L6MUX21 i1580 (.D0(n1761), .D1(n1762), .SD(address[2]), .Z(n1766));
    L6MUX21 i1484 (.D0(n1662), .D1(n1663), .SD(address[2]), .Z(n1670));
    L6MUX21 i1579 (.D0(n1759), .D1(n1760), .SD(address[2]), .Z(n1765));
    L6MUX21 i1578 (.D0(n1757), .D1(n1758), .SD(address[2]), .Z(n1764));
    L6MUX21 i1577 (.D0(n1755), .D1(n1756), .SD(address[2]), .Z(n1763));
    L6MUX21 i1270 (.D0(n1451), .D1(n1452), .SD(address[2]), .Z(n1456));
    L6MUX21 i1269 (.D0(n1449), .D1(n1450), .SD(address[2]), .Z(n1455));
    L6MUX21 i1268 (.D0(n1447), .D1(n1448), .SD(address[2]), .Z(n1454));
    L6MUX21 i1267 (.D0(n1445), .D1(n1446), .SD(address[2]), .Z(n1453));
    L6MUX21 i1239 (.D0(n1420), .D1(n1421), .SD(address[2]), .Z(n1425));
    L6MUX21 i1238 (.D0(n1418), .D1(n1419), .SD(address[2]), .Z(n1424));
    L6MUX21 i1237 (.D0(n1416), .D1(n1417), .SD(address[2]), .Z(n1423));
    L6MUX21 i1236 (.D0(n1414), .D1(n1415), .SD(address[2]), .Z(n1422));
    L6MUX21 i1456 (.D0(n1637), .D1(n1638), .SD(address[2]), .Z(n1642));
    L6MUX21 i1455 (.D0(n1635), .D1(n1636), .SD(address[2]), .Z(n1641));
    L6MUX21 i1454 (.D0(n1633), .D1(n1634), .SD(address[2]), .Z(n1640));
    L6MUX21 i1453 (.D0(n1631), .D1(n1632), .SD(address[2]), .Z(n1639));
    L6MUX21 i1208 (.D0(n1389), .D1(n1390), .SD(address[2]), .Z(n1394));
    L6MUX21 i1207 (.D0(n1387), .D1(n1388), .SD(address[2]), .Z(n1393));
    L6MUX21 i1206 (.D0(n1385), .D1(n1386), .SD(address[2]), .Z(n1392));
    L6MUX21 i1205 (.D0(n1383), .D1(n1384), .SD(address[2]), .Z(n1391));
    L6MUX21 i1425 (.D0(n1606), .D1(n1607), .SD(address[2]), .Z(n1611));
    L6MUX21 i1424 (.D0(n1604), .D1(n1605), .SD(address[2]), .Z(n1610));
    L6MUX21 i1549 (.D0(n1730), .D1(n1731), .SD(address[2]), .Z(n1735));
    L6MUX21 i1423 (.D0(n1602), .D1(n1603), .SD(address[2]), .Z(n1609));
    L6MUX21 i1422 (.D0(n1600), .D1(n1601), .SD(address[2]), .Z(n1608));
    L6MUX21 i1548 (.D0(n1728), .D1(n1729), .SD(address[2]), .Z(n1734));
    L6MUX21 i1547 (.D0(n1726), .D1(n1727), .SD(address[2]), .Z(n1733));
    L6MUX21 i1177 (.D0(n1358), .D1(n1359), .SD(address[2]), .Z(n1363));
    L6MUX21 i1176 (.D0(n1356), .D1(n1357), .SD(address[2]), .Z(n1362));
    L6MUX21 i1175 (.D0(n1354), .D1(n1355), .SD(address[2]), .Z(n1361));
    L6MUX21 i1546 (.D0(n1724), .D1(n1725), .SD(address[2]), .Z(n1732));
    L6MUX21 i1174 (.D0(n1352), .D1(n1353), .SD(address[2]), .Z(n1360));
    L6MUX21 i1611 (.D0(n1792), .D1(n1793), .SD(address[2]), .Z(n1797));
    L6MUX21 i1643 (.D0(n1825), .D1(n1826), .SD(address[3]), .Z(n1829));
    L6MUX21 i1396 (.D0(n1579), .D1(n1580), .SD(address[3]), .Z(n1582));
    L6MUX21 i1395 (.D0(n1577), .D1(n1578), .SD(address[3]), .Z(n1581));
    L6MUX21 i1365 (.D0(n1548), .D1(n1549), .SD(address[3]), .Z(n1551));
    L6MUX21 i1364 (.D0(n1546), .D1(n1547), .SD(address[3]), .Z(n1550));
    L6MUX21 i1520 (.D0(n1703), .D1(n1704), .SD(address[3]), .Z(n1706));
    L6MUX21 i1519 (.D0(n1701), .D1(n1702), .SD(address[3]), .Z(n1705));
    L6MUX21 i1334 (.D0(n1517), .D1(n1518), .SD(address[3]), .Z(n1520));
    L6MUX21 i1333 (.D0(n1515), .D1(n1516), .SD(address[3]), .Z(n1519));
    L6MUX21 i1582 (.D0(n1765), .D1(n1766), .SD(address[3]), .Z(n1768));
    L6MUX21 i1303 (.D0(n1486), .D1(n1487), .SD(address[3]), .Z(n1489));
    L6MUX21 i1302 (.D0(n1484), .D1(n1485), .SD(address[3]), .Z(n1488));
    L6MUX21 i1489 (.D0(n1672), .D1(n1673), .SD(address[3]), .Z(n1675));
    L6MUX21 i1488 (.D0(n1670), .D1(n1671), .SD(address[3]), .Z(n1674));
    L6MUX21 i1581 (.D0(n1763), .D1(n1764), .SD(address[3]), .Z(n1767));
    L6MUX21 i1272 (.D0(n1455), .D1(n1456), .SD(address[3]), .Z(n1458));
    L6MUX21 i1271 (.D0(n1453), .D1(n1454), .SD(address[3]), .Z(n1457));
    L6MUX21 i1241 (.D0(n1424), .D1(n1425), .SD(address[3]), .Z(n1427));
    L6MUX21 i1240 (.D0(n1422), .D1(n1423), .SD(address[3]), .Z(n1426));
    L6MUX21 i1458 (.D0(n1641), .D1(n1642), .SD(address[3]), .Z(n1644));
    L6MUX21 i1457 (.D0(n1639), .D1(n1640), .SD(address[3]), .Z(n1643));
    L6MUX21 i1210 (.D0(n1393), .D1(n1394), .SD(address[3]), .Z(n1396));
    L6MUX21 i1209 (.D0(n1391), .D1(n1392), .SD(address[3]), .Z(n1395));
    L6MUX21 i1551 (.D0(n1734), .D1(n1735), .SD(address[3]), .Z(n1737));
    L6MUX21 i1427 (.D0(n1610), .D1(n1611), .SD(address[3]), .Z(n1613));
    L6MUX21 i1426 (.D0(n1608), .D1(n1609), .SD(address[3]), .Z(n1612));
    L6MUX21 i1550 (.D0(n1732), .D1(n1733), .SD(address[3]), .Z(n1736));
    L6MUX21 i1613 (.D0(n1796), .D1(n1797), .SD(address[3]), .Z(n1799));
    L6MUX21 i1179 (.D0(n1362), .D1(n1363), .SD(address[3]), .Z(n1365));
    L6MUX21 i1612 (.D0(n1794), .D1(n1795), .SD(address[3]), .Z(n1798));
    L6MUX21 i1178 (.D0(n1360), .D1(n1361), .SD(address[3]), .Z(n1364));
    L6MUX21 i1644 (.D0(n1827), .D1(n1828), .SD(address[3]), .Z(n1830));
    PFUMX i94611_i1 (.BLUT(n1366), .ALUT(n1831), .C0(address[5]), .Z(data_7__N_84[7]));
    PFUMX i95214_i1 (.BLUT(n1397), .ALUT(n1800), .C0(address[5]), .Z(data_7__N_84[2]));
    PFUMX i95817_i1 (.BLUT(n1428), .ALUT(n1769), .C0(address[5]), .Z(data_7__N_84[6]));
    PFUMX i96420_i1 (.BLUT(n1459), .ALUT(n1738), .C0(address[5]), .Z(data_7__N_84[5]));
    PFUMX i97023_i1 (.BLUT(n1490), .ALUT(n1707), .C0(address[5]), .Z(data_7__N_84[4]));
    PFUMX i97626_i1 (.BLUT(n1521), .ALUT(n1676), .C0(address[5]), .Z(data_7__N_84[3]));
    PFUMX i98229_i1 (.BLUT(n1552), .ALUT(n1645), .C0(address[5]), .Z(data_7__N_84[0]));
    PFUMX i98832_i1 (.BLUT(n1583), .ALUT(n1614), .C0(address[5]), .Z(data_7__N_84[1]));
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module CPU8BIT2
//

module CPU8BIT2 (address, clk_c, akku_o_c_0, n1916, data, akku_o_c_7, 
            akku_o_c_6, akku_o_c_5, akku_o_c_4, \states_2__N_71[2] , 
            akku_o_c_3, akku_o_c_2, akku_o_c_1, reset_c, data_7__N_97, 
            n1895, n1905, n1328, n1898, mem_0__7__N_101, n1899, 
            mem_15__7__N_148, n1302, mem_12__7__N_139, mem_7__7__N_124, 
            n1906, mem_56__7__N_271, n1327, mem_58__7__N_277, mem_59__7__N_280, 
            mem_60__7__N_283, mem_63__7__N_292, n1902, mem_48__7__N_247, 
            mem_50__7__N_253, mem_51__7__N_256, mem_52__7__N_259, mem_55__7__N_268, 
            n1901, mem_40__7__N_223, mem_42__7__N_229, mem_43__7__N_232, 
            mem_44__7__N_235, mem_47__7__N_244, n1911, mem_32__7__N_199, 
            mem_34__7__N_205, mem_35__7__N_208, mem_36__7__N_211, mem_39__7__N_220, 
            n1910, mem_24__7__N_175, mem_26__7__N_181, mem_27__7__N_184, 
            akku_o_c_8, mem_28__7__N_187, \states_2__N_71[0] , n1896, 
            mem_31__7__N_196, n1900, mem_16__7__N_151, mem_18__7__N_157, 
            mem_19__7__N_160, mem_20__7__N_163, mem_23__7__N_172, mem_8__7__N_127, 
            mem_10__7__N_133, mem_11__7__N_136, mem_4__7__N_115, mem_3__7__N_112, 
            mem_2__7__N_109, GND_net);
    output [5:0]address;
    input clk_c;
    output akku_o_c_0;
    input n1916;
    input [7:0]data;
    output akku_o_c_7;
    output akku_o_c_6;
    output akku_o_c_5;
    output akku_o_c_4;
    input \states_2__N_71[2] ;
    output akku_o_c_3;
    output akku_o_c_2;
    output akku_o_c_1;
    input reset_c;
    output data_7__N_97;
    input n1895;
    output n1905;
    input n1328;
    input n1898;
    output mem_0__7__N_101;
    input n1899;
    output mem_15__7__N_148;
    input n1302;
    output mem_12__7__N_139;
    output mem_7__7__N_124;
    input n1906;
    output mem_56__7__N_271;
    input n1327;
    output mem_58__7__N_277;
    output mem_59__7__N_280;
    output mem_60__7__N_283;
    output mem_63__7__N_292;
    input n1902;
    output mem_48__7__N_247;
    output mem_50__7__N_253;
    output mem_51__7__N_256;
    output mem_52__7__N_259;
    output mem_55__7__N_268;
    input n1901;
    output mem_40__7__N_223;
    output mem_42__7__N_229;
    output mem_43__7__N_232;
    output mem_44__7__N_235;
    output mem_47__7__N_244;
    input n1911;
    output mem_32__7__N_199;
    output mem_34__7__N_205;
    output mem_35__7__N_208;
    output mem_36__7__N_211;
    output mem_39__7__N_220;
    input n1910;
    output mem_24__7__N_175;
    output mem_26__7__N_181;
    output mem_27__7__N_184;
    output akku_o_c_8;
    output mem_28__7__N_187;
    input \states_2__N_71[0] ;
    output n1896;
    output mem_31__7__N_196;
    input n1900;
    output mem_16__7__N_151;
    output mem_18__7__N_157;
    output mem_19__7__N_160;
    output mem_20__7__N_163;
    output mem_23__7__N_172;
    output mem_8__7__N_127;
    output mem_10__7__N_133;
    output mem_11__7__N_136;
    output mem_4__7__N_115;
    output mem_3__7__N_112;
    output mem_2__7__N_109;
    input GND_net;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(8[13:16])
    wire mem_0__7__N_101 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_0__7__N_101 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_15__7__N_148 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_15__7__N_148 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_12__7__N_139 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_12__7__N_139 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_7__7__N_124 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_7__7__N_124 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_56__7__N_271 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_56__7__N_271 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_58__7__N_277 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_58__7__N_277 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_59__7__N_280 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_59__7__N_280 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_60__7__N_283 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_60__7__N_283 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_63__7__N_292 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_63__7__N_292 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_48__7__N_247 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_48__7__N_247 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_50__7__N_253 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_50__7__N_253 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_51__7__N_256 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_51__7__N_256 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_52__7__N_259 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_52__7__N_259 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_55__7__N_268 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_55__7__N_268 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_40__7__N_223 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_40__7__N_223 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_42__7__N_229 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_42__7__N_229 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_43__7__N_232 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_43__7__N_232 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_44__7__N_235 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_44__7__N_235 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_47__7__N_244 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_47__7__N_244 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_32__7__N_199 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_32__7__N_199 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_34__7__N_205 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_34__7__N_205 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_35__7__N_208 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_35__7__N_208 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_36__7__N_211 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_36__7__N_211 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_39__7__N_220 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_39__7__N_220 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_24__7__N_175 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_24__7__N_175 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_26__7__N_181 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_26__7__N_181 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_27__7__N_184 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_27__7__N_184 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_28__7__N_187 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_28__7__N_187 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_31__7__N_196 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_31__7__N_196 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_16__7__N_151 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_16__7__N_151 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_18__7__N_157 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_18__7__N_157 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_19__7__N_160 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_19__7__N_160 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_20__7__N_163 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_20__7__N_163 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_23__7__N_172 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_23__7__N_172 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_8__7__N_127 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_8__7__N_127 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_10__7__N_133 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_10__7__N_133 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_11__7__N_136 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_11__7__N_136 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_4__7__N_115 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_4__7__N_115 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_3__7__N_112 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_3__7__N_112 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_2__7__N_109 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_2__7__N_109 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [5:0]adress_5__N_3;
    
    wire clk_c_enable_15;
    wire [8:0]n198;
    wire [5:0]pc;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(23[15:17])
    
    wire clk_c_enable_7;
    wire [2:0]states;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(25[15:21])
    wire [8:0]n228;
    
    wire n1908, n605;
    wire [2:0]n297;
    wire [5:0]pc_5__N_30;
    
    wire n1999, n1913, n1903, n1917, n876, clk_c_enable_8, n572, 
        n588, n570, n592, n590, n1907, n1281, n1280, n1279, 
        n1278, n1277;
    
    FD1S3AX adreg_i0 (.D(adress_5__N_3[0]), .CK(clk_c), .Q(address[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam adreg_i0.GSR = "ENABLED";
    FD1P3AX akku_i0_i1 (.D(n198[0]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_0)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam akku_i0_i1.GSR = "ENABLED";
    FD1P3AX pc_i0_i0 (.D(n1916), .SP(clk_c_enable_7), .CK(clk_c), .Q(pc[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam pc_i0_i0.GSR = "ENABLED";
    LUT4 mux_105_i1_4_lut_4_lut (.A(states[0]), .B(data[0]), .C(akku_o_c_0), 
         .D(n228[0]), .Z(n198[0])) /* synthesis lut_function=(!(A (B+(C))+!A !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[33:48])
    defparam mux_105_i1_4_lut_4_lut.init = 16'h5702;
    LUT4 mux_105_i8_4_lut_4_lut (.A(states[0]), .B(data[7]), .C(akku_o_c_7), 
         .D(n228[7]), .Z(n198[7])) /* synthesis lut_function=(!(A (B+(C))+!A !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[33:48])
    defparam mux_105_i8_4_lut_4_lut.init = 16'h5702;
    LUT4 mux_105_i7_4_lut_4_lut (.A(states[0]), .B(data[6]), .C(akku_o_c_6), 
         .D(n228[6]), .Z(n198[6])) /* synthesis lut_function=(!(A (B+(C))+!A !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[33:48])
    defparam mux_105_i7_4_lut_4_lut.init = 16'h5702;
    LUT4 mux_105_i6_4_lut_4_lut (.A(states[0]), .B(data[5]), .C(akku_o_c_5), 
         .D(n228[5]), .Z(n198[5])) /* synthesis lut_function=(!(A (B+(C))+!A !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[33:48])
    defparam mux_105_i6_4_lut_4_lut.init = 16'h5702;
    LUT4 mux_105_i5_4_lut_4_lut (.A(states[0]), .B(data[4]), .C(akku_o_c_4), 
         .D(n228[4]), .Z(n198[4])) /* synthesis lut_function=(!(A (B+(C))+!A !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[33:48])
    defparam mux_105_i5_4_lut_4_lut.init = 16'h5702;
    FD1S3IX states__i2 (.D(\states_2__N_71[2] ), .CK(clk_c), .CD(n1908), 
            .Q(states[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam states__i2.GSR = "ENABLED";
    FD1S3IX states__i1 (.D(n297[1]), .CK(clk_c), .CD(n605), .Q(states[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam states__i1.GSR = "ENABLED";
    LUT4 mux_105_i4_4_lut_4_lut (.A(states[0]), .B(data[3]), .C(akku_o_c_3), 
         .D(n228[3]), .Z(n198[3])) /* synthesis lut_function=(!(A (B+(C))+!A !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[33:48])
    defparam mux_105_i4_4_lut_4_lut.init = 16'h5702;
    LUT4 mux_105_i3_4_lut_4_lut (.A(states[0]), .B(data[2]), .C(akku_o_c_2), 
         .D(n228[2]), .Z(n198[2])) /* synthesis lut_function=(!(A (B+(C))+!A !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[33:48])
    defparam mux_105_i3_4_lut_4_lut.init = 16'h5702;
    LUT4 mux_105_i2_4_lut_4_lut (.A(states[0]), .B(data[1]), .C(akku_o_c_1), 
         .D(n228[1]), .Z(n198[1])) /* synthesis lut_function=(!(A (B+(C))+!A !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[33:48])
    defparam mux_105_i2_4_lut_4_lut.init = 16'h5702;
    FD1P3AX pc_i0_i5 (.D(pc_5__N_30[5]), .SP(clk_c_enable_7), .CK(clk_c), 
            .Q(pc[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam pc_i0_i5.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_87 (.A(reset_c), .B(clk_c), .Z(n1999)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_rep_87.init = 16'h2222;
    LUT4 i1_3_lut_3_lut_2_lut_3_lut_4_lut (.A(reset_c), .B(clk_c), .C(states[0]), 
         .D(states[1]), .Z(data_7__N_97)) /* synthesis lut_function=(!((B+!((D)+!C))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_3_lut_3_lut_2_lut_3_lut_4_lut.init = 16'h2202;
    LUT4 i191_2_lut_3_lut_4_lut (.A(address[2]), .B(n1913), .C(address[4]), 
         .D(address[3]), .Z(pc_5__N_30[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i191_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i1_3_lut_4_lut (.A(data[6]), .B(n1895), .C(n1908), .D(data[5]), 
         .Z(n605)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (C)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(37[13:17])
    defparam i1_3_lut_4_lut.init = 16'hf0f8;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n1905), .B(n1999), .C(n1328), .D(n1898), 
         .Z(mem_0__7__N_101)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i13_3_lut (.A(states[1]), .B(states[0]), .C(states[2]), .Z(clk_c_enable_15)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam i13_3_lut.init = 16'h3a3a;
    LUT4 i1_2_lut_3_lut_4_lut_adj_8 (.A(n1905), .B(n1999), .C(n1903), 
         .D(n1899), .Z(mem_15__7__N_148)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_8.init = 16'h0040;
    LUT4 i198_3_lut_4_lut (.A(address[3]), .B(n1903), .C(address[4]), 
         .D(address[5]), .Z(pc_5__N_30[5])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i198_3_lut_4_lut.init = 16'h7f80;
    LUT4 pc_5__I_0_100_i6_3_lut_4_lut (.A(states[1]), .B(n1917), .C(pc[5]), 
         .D(data[5]), .Z(adress_5__N_3[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[33:48])
    defparam pc_5__I_0_100_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pc_5__I_0_100_i4_3_lut_4_lut (.A(states[1]), .B(n1917), .C(pc[3]), 
         .D(data[3]), .Z(adress_5__N_3[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[33:48])
    defparam pc_5__I_0_100_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pc_5__I_0_100_i5_3_lut_4_lut (.A(states[1]), .B(n1917), .C(pc[4]), 
         .D(data[4]), .Z(adress_5__N_3[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[33:48])
    defparam pc_5__I_0_100_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pc_5__I_0_100_i1_3_lut_4_lut (.A(states[1]), .B(n1917), .C(pc[0]), 
         .D(data[0]), .Z(adress_5__N_3[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[33:48])
    defparam pc_5__I_0_100_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pc_5__I_0_100_i3_3_lut_4_lut (.A(states[1]), .B(n1917), .C(pc[2]), 
         .D(data[2]), .Z(adress_5__N_3[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[33:48])
    defparam pc_5__I_0_100_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_9 (.A(n1905), .B(n1999), .C(n1302), 
         .D(n1899), .Z(mem_12__7__N_139)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_9.init = 16'h0004;
    LUT4 pc_5__I_0_100_i2_3_lut_4_lut (.A(states[1]), .B(n1917), .C(pc[1]), 
         .D(data[1]), .Z(adress_5__N_3[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[33:48])
    defparam pc_5__I_0_100_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_10 (.A(n1905), .B(n1999), .C(n1903), 
         .D(n1898), .Z(mem_7__7__N_124)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_10.init = 16'h0040;
    LUT4 i1_2_lut_3_lut_4_lut_adj_11 (.A(n1905), .B(n1999), .C(n1328), 
         .D(n1906), .Z(mem_56__7__N_271)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_11.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_12 (.A(n1905), .B(n1999), .C(n1327), 
         .D(n1906), .Z(mem_58__7__N_277)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_12.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_13 (.A(n1905), .B(n1999), .C(n876), 
         .D(n1906), .Z(mem_59__7__N_280)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_13.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_14 (.A(n1905), .B(n1999), .C(n1302), 
         .D(n1906), .Z(mem_60__7__N_283)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_14.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_15 (.A(n1905), .B(n1999), .C(n1903), 
         .D(n1906), .Z(mem_63__7__N_292)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_15.init = 16'h4000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_16 (.A(n1905), .B(n1999), .C(n1328), 
         .D(n1902), .Z(mem_48__7__N_247)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_16.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_17 (.A(n1905), .B(n1999), .C(n1327), 
         .D(n1902), .Z(mem_50__7__N_253)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_17.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_18 (.A(n1905), .B(n1999), .C(n876), 
         .D(n1902), .Z(mem_51__7__N_256)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_18.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_19 (.A(n1905), .B(n1999), .C(n1302), 
         .D(n1902), .Z(mem_52__7__N_259)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_19.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_20 (.A(n1905), .B(n1999), .C(n1903), 
         .D(n1902), .Z(mem_55__7__N_268)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_20.init = 16'h0040;
    LUT4 i1_2_lut_3_lut_4_lut_adj_21 (.A(n1905), .B(n1999), .C(n1328), 
         .D(n1901), .Z(mem_40__7__N_223)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_21.init = 16'h0004;
    LUT4 i172_2_lut_rep_82 (.A(address[1]), .B(address[0]), .Z(n1913)) /* synthesis lut_function=(A (B)) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i172_2_lut_rep_82.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_22 (.A(n1905), .B(n1999), .C(n1327), 
         .D(n1901), .Z(mem_42__7__N_229)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_22.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_23 (.A(n1905), .B(n1999), .C(n876), 
         .D(n1901), .Z(mem_43__7__N_232)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_23.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_24 (.A(n1905), .B(n1999), .C(n1302), 
         .D(n1901), .Z(mem_44__7__N_235)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_24.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_25 (.A(n1905), .B(n1999), .C(n1903), 
         .D(n1901), .Z(mem_47__7__N_244)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_25.init = 16'h0040;
    LUT4 i179_2_lut_rep_72_3_lut (.A(address[1]), .B(address[0]), .C(address[2]), 
         .Z(n1903)) /* synthesis lut_function=(A (B (C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i179_2_lut_rep_72_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_26 (.A(n1905), .B(n1999), .C(n1328), 
         .D(n1911), .Z(mem_32__7__N_199)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_26.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_27 (.A(n1905), .B(n1999), .C(n1327), 
         .D(n1911), .Z(mem_34__7__N_205)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_27.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_28 (.A(n1905), .B(n1999), .C(n876), 
         .D(n1911), .Z(mem_35__7__N_208)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_28.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_29 (.A(n1905), .B(n1999), .C(n1302), 
         .D(n1911), .Z(mem_36__7__N_211)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_29.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_30 (.A(n1905), .B(n1999), .C(n1903), 
         .D(n1911), .Z(mem_39__7__N_220)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_30.init = 16'h0040;
    LUT4 i1_2_lut_3_lut_4_lut_adj_31 (.A(n1905), .B(n1999), .C(n1328), 
         .D(n1910), .Z(mem_24__7__N_175)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_31.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_32 (.A(n1905), .B(n1999), .C(n1327), 
         .D(n1910), .Z(mem_26__7__N_181)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_32.init = 16'h0004;
    LUT4 i1_2_lut_3_lut (.A(address[1]), .B(address[0]), .C(address[2]), 
         .Z(n876)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i1_2_lut_3_lut.init = 16'hf7f7;
    FD1P3AX pc_i0_i4 (.D(pc_5__N_30[4]), .SP(clk_c_enable_7), .CK(clk_c), 
            .Q(pc[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam pc_i0_i4.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_33 (.A(n1905), .B(n1999), .C(n876), 
         .D(n1910), .Z(mem_27__7__N_184)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_33.init = 16'h0004;
    FD1P3AX pc_i0_i3 (.D(pc_5__N_30[3]), .SP(clk_c_enable_7), .CK(clk_c), 
            .Q(pc[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam pc_i0_i3.GSR = "ENABLED";
    FD1P3AX pc_i0_i2 (.D(pc_5__N_30[2]), .SP(clk_c_enable_7), .CK(clk_c), 
            .Q(pc[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam pc_i0_i2.GSR = "ENABLED";
    FD1P3AX pc_i0_i1 (.D(pc_5__N_30[1]), .SP(clk_c_enable_7), .CK(clk_c), 
            .Q(pc[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam pc_i0_i1.GSR = "ENABLED";
    FD1P3AX akku_i0_i9 (.D(n198[8]), .SP(clk_c_enable_8), .CK(clk_c), 
            .Q(akku_o_c_8)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam akku_i0_i9.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_34 (.A(n1905), .B(n1999), .C(n1302), 
         .D(n1910), .Z(mem_28__7__N_187)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_34.init = 16'h0004;
    FD1S3IX states__i0 (.D(\states_2__N_71[0] ), .CK(clk_c), .CD(n1908), 
            .Q(states[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam states__i0.GSR = "ENABLED";
    FD1P3AX akku_i0_i8 (.D(n198[7]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_7)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam akku_i0_i8.GSR = "ENABLED";
    FD1P3AX akku_i0_i7 (.D(n198[6]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_6)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam akku_i0_i7.GSR = "ENABLED";
    FD1P3AX akku_i0_i6 (.D(n198[5]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_5)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam akku_i0_i6.GSR = "ENABLED";
    FD1P3AX akku_i0_i5 (.D(n198[4]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_4)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam akku_i0_i5.GSR = "ENABLED";
    FD1P3AX akku_i0_i4 (.D(n198[3]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_3)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam akku_i0_i4.GSR = "ENABLED";
    FD1P3AX akku_i0_i3 (.D(n198[2]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_2)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam akku_i0_i3.GSR = "ENABLED";
    FD1P3AX akku_i0_i2 (.D(n198[1]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(akku_o_c_1)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam akku_i0_i2.GSR = "ENABLED";
    FD1S3AX adreg_i5 (.D(adress_5__N_3[5]), .CK(clk_c), .Q(address[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam adreg_i5.GSR = "ENABLED";
    FD1S3AX adreg_i4 (.D(adress_5__N_3[4]), .CK(clk_c), .Q(address[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam adreg_i4.GSR = "ENABLED";
    LUT4 i177_2_lut_3_lut (.A(address[1]), .B(address[0]), .C(address[2]), 
         .Z(pc_5__N_30[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i177_2_lut_3_lut.init = 16'h7878;
    LUT4 i184_2_lut_3_lut_4_lut (.A(address[1]), .B(address[0]), .C(address[3]), 
         .D(address[2]), .Z(pc_5__N_30[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i184_2_lut_3_lut_4_lut.init = 16'h78f0;
    FD1S3AX adreg_i3 (.D(adress_5__N_3[3]), .CK(clk_c), .Q(address[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam adreg_i3.GSR = "ENABLED";
    FD1S3AX adreg_i2 (.D(adress_5__N_3[2]), .CK(clk_c), .Q(address[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam adreg_i2.GSR = "ENABLED";
    FD1S3AX adreg_i1 (.D(adress_5__N_3[1]), .CK(clk_c), .Q(address[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(29[9] 79[16])
    defparam adreg_i1.GSR = "ENABLED";
    LUT4 i1_3_lut (.A(data[5]), .B(data[7]), .C(data[6]), .Z(n297[1])) /* synthesis lut_function=(A ((C)+!B)+!A !(B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(37[13:17])
    defparam i1_3_lut.init = 16'hb3b3;
    LUT4 i1_2_lut_rep_65_3_lut_4_lut (.A(states[1]), .B(states[0]), .C(n1999), 
         .D(states[2]), .Z(n1896)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(86[65:80])
    defparam i1_2_lut_rep_65_3_lut_4_lut.init = 16'h0040;
    LUT4 i170_2_lut (.A(address[1]), .B(address[0]), .Z(pc_5__N_30[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i170_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_rep_74_3_lut (.A(states[1]), .B(states[0]), .C(states[2]), 
         .Z(n1905)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(86[65:80])
    defparam i1_2_lut_rep_74_3_lut.init = 16'hfbfb;
    LUT4 i1_2_lut (.A(address[4]), .B(states[1]), .Z(n572)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_adj_35 (.A(address[2]), .B(states[1]), .Z(n588)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_35.init = 16'h6666;
    LUT4 i1_2_lut_adj_36 (.A(address[3]), .B(states[1]), .Z(n570)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_36.init = 16'h6666;
    LUT4 i1_2_lut_adj_37 (.A(address[0]), .B(states[1]), .Z(n592)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_37.init = 16'h6666;
    LUT4 i1_2_lut_adj_38 (.A(address[1]), .B(states[1]), .Z(n590)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_38.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut_adj_39 (.A(n1905), .B(n1999), .C(n1903), 
         .D(n1910), .Z(mem_31__7__N_196)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_39.init = 16'h0040;
    LUT4 i1_2_lut_3_lut_4_lut_adj_40 (.A(n1905), .B(n1999), .C(n1328), 
         .D(n1900), .Z(mem_16__7__N_151)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_40.init = 16'h0004;
    LUT4 i1_2_lut_rep_86 (.A(states[2]), .B(states[0]), .Z(n1917)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[33:48])
    defparam i1_2_lut_rep_86.init = 16'heeee;
    LUT4 i113_2_lut_rep_76_3_lut (.A(states[2]), .B(states[0]), .C(states[1]), 
         .Z(n1907)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[33:48])
    defparam i113_2_lut_rep_76_3_lut.init = 16'h1010;
    LUT4 i19_4_lut_4_lut_4_lut_3_lut (.A(states[2]), .B(states[0]), .C(states[1]), 
         .Z(clk_c_enable_8)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[33:48])
    defparam i19_4_lut_4_lut_4_lut_3_lut.init = 16'h3a3a;
    LUT4 i1_2_lut_3_lut_4_lut_adj_41 (.A(n1905), .B(n1999), .C(n1327), 
         .D(n1900), .Z(mem_18__7__N_157)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_41.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_42 (.A(n1905), .B(n1999), .C(n876), 
         .D(n1900), .Z(mem_19__7__N_160)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_42.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_43 (.A(n1905), .B(n1999), .C(n1302), 
         .D(n1900), .Z(mem_20__7__N_163)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_43.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_44 (.A(n1905), .B(n1999), .C(n1903), 
         .D(n1900), .Z(mem_23__7__N_172)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_44.init = 16'h0040;
    LUT4 i1_2_lut_3_lut_4_lut_2_lut (.A(states[0]), .B(n228[8]), .Z(n198[8])) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[33:48])
    defparam i1_2_lut_3_lut_4_lut_2_lut.init = 16'h4444;
    LUT4 i2_2_lut_rep_77_3_lut (.A(states[2]), .B(states[0]), .C(states[1]), 
         .Z(n1908)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[33:48])
    defparam i2_2_lut_rep_77_3_lut.init = 16'hfefe;
    LUT4 i736_1_lut_2_lut_3_lut (.A(states[2]), .B(states[0]), .C(states[1]), 
         .Z(clk_c_enable_7)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[33:48])
    defparam i736_1_lut_2_lut_3_lut.init = 16'h0101;
    LUT4 i1_2_lut_3_lut_4_lut_adj_45 (.A(n1905), .B(n1999), .C(n1328), 
         .D(n1899), .Z(mem_8__7__N_127)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_45.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_46 (.A(n1905), .B(n1999), .C(n1327), 
         .D(n1899), .Z(mem_10__7__N_133)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_46.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_47 (.A(n1905), .B(n1999), .C(n876), 
         .D(n1899), .Z(mem_11__7__N_136)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_47.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_48 (.A(n1905), .B(n1999), .C(n1302), 
         .D(n1898), .Z(mem_4__7__N_115)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_48.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_49 (.A(n1905), .B(n1999), .C(n876), 
         .D(n1898), .Z(mem_3__7__N_112)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_49.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_50 (.A(n1905), .B(n1999), .C(n1327), 
         .D(n1898), .Z(mem_2__7__N_109)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(87[21:60])
    defparam i1_2_lut_3_lut_4_lut_adj_50.init = 16'h0004;
    CCU2D add_132_11 (.A0(n1917), .B0(states[1]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n1281), 
          .S0(n228[8]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[13] 53[22])
    defparam add_132_11.INIT0 = 16'h7888;
    defparam add_132_11.INIT1 = 16'h0000;
    defparam add_132_11.INJECT1_0 = "NO";
    defparam add_132_11.INJECT1_1 = "NO";
    CCU2D add_132_9 (.A0(akku_o_c_6), .B0(data[6]), .C0(n1917), .D0(states[1]), 
          .A1(akku_o_c_7), .B1(data[7]), .C1(n1917), .D1(states[1]), 
          .CIN(n1280), .COUT(n1281), .S0(n228[6]), .S1(n228[7]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[13] 53[22])
    defparam add_132_9.INIT0 = 16'h56aa;
    defparam add_132_9.INIT1 = 16'h56aa;
    defparam add_132_9.INJECT1_0 = "NO";
    defparam add_132_9.INJECT1_1 = "NO";
    CCU2D add_132_7 (.A0(akku_o_c_4), .B0(n1907), .C0(data[4]), .D0(n572), 
          .A1(akku_o_c_5), .B1(data[5]), .C1(n1917), .D1(states[1]), 
          .CIN(n1279), .COUT(n1280), .S0(n228[4]), .S1(n228[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[13] 53[22])
    defparam add_132_7.INIT0 = 16'h596a;
    defparam add_132_7.INIT1 = 16'h56aa;
    defparam add_132_7.INJECT1_0 = "NO";
    defparam add_132_7.INJECT1_1 = "NO";
    CCU2D add_132_5 (.A0(akku_o_c_2), .B0(n1907), .C0(data[2]), .D0(n588), 
          .A1(akku_o_c_3), .B1(n1907), .C1(data[3]), .D1(n570), .CIN(n1278), 
          .COUT(n1279), .S0(n228[2]), .S1(n228[3]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[13] 53[22])
    defparam add_132_5.INIT0 = 16'h596a;
    defparam add_132_5.INIT1 = 16'h596a;
    defparam add_132_5.INJECT1_0 = "NO";
    defparam add_132_5.INJECT1_1 = "NO";
    CCU2D add_132_3 (.A0(akku_o_c_0), .B0(n1907), .C0(data[0]), .D0(n592), 
          .A1(akku_o_c_1), .B1(n1907), .C1(data[1]), .D1(n590), .CIN(n1277), 
          .COUT(n1278), .S0(n228[0]), .S1(n228[1]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[13] 53[22])
    defparam add_132_3.INIT0 = 16'h596a;
    defparam add_132_3.INIT1 = 16'h596a;
    defparam add_132_3.INJECT1_0 = "NO";
    defparam add_132_3.INJECT1_1 = "NO";
    CCU2D add_132_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1917), .B1(states[1]), .C1(GND_net), .D1(GND_net), .COUT(n1277));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[13] 53[22])
    defparam add_132_1.INIT0 = 16'hF000;
    defparam add_132_1.INIT1 = 16'h7777;
    defparam add_132_1.INJECT1_0 = "NO";
    defparam add_132_1.INJECT1_1 = "NO";
    
endmodule
