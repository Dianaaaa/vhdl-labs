// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.11.0.396.4
// Netlist written on Mon Nov 23 13:57:24 2020
//
// Verilog Description of module cpu2system
//

module cpu2system (clk, reset, akku_o);   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(7[8:18])
    input clk;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(8[13:16])
    input reset;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(9[13:18])
    output [8:0]akku_o;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(8[13:16])
    
    wire GND_net, VCC_net, reset_c, akku_o_c_8, akku_o_c_7, akku_o_c_6, 
        akku_o_c_5, akku_o_c_4, akku_o_c_3, akku_o_c_2, akku_o_c_1, 
        akku_o_c_0;
    wire [7:0]data;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(37[13:17])
    wire [2:0]states;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(22[15:21])
    wire [5:0]address;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(24[9:16])
    wire [7:0]data_7__N_89;
    
    wire data_7__N_102, n46237, n46211, n23757;
    
    VHI i33735 (.Z(VCC_net));
    IB reset_pad (.I(reset), .O(reset_c));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(9[13:18])
    IB clk_pad (.I(clk), .O(clk_c));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(8[13:16])
    OB akku_o_pad_0 (.I(akku_o_c_0), .O(akku_o[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_1 (.I(akku_o_c_1), .O(akku_o[1]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_2 (.I(akku_o_c_2), .O(akku_o[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_3 (.I(akku_o_c_3), .O(akku_o[3]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_4 (.I(akku_o_c_4), .O(akku_o[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_5 (.I(akku_o_c_5), .O(akku_o[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_6 (.I(akku_o_c_6), .O(akku_o[6]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_7 (.I(akku_o_c_7), .O(akku_o[7]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    OB akku_o_pad_8 (.I(akku_o_c_8), .O(akku_o[8]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    VLO i1 (.Z(GND_net));
    GSR GSR_INST (.GSR(reset_c));
    TSALL TSALL_INST (.TSALL(GND_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    CPU8BIT2 CPU (.states({Open_0, Open_1, states[0]}), .clk_c(clk_c), 
            .akku_o_c_0(akku_o_c_0), .address({address}), .data({data}), 
            .GND_net(GND_net), .akku_o_c_4(akku_o_c_4), .akku_o_c_1(akku_o_c_1), 
            .akku_o_c_2(akku_o_c_2), .akku_o_c_3(akku_o_c_3), .\states[1] (states[1]), 
            .akku_o_c_7(akku_o_c_7), .data_7__N_89({data_7__N_89}), .data_7__N_102(data_7__N_102), 
            .akku_o_c_5(akku_o_c_5), .akku_o_c_6(akku_o_c_6), .VCC_net(VCC_net), 
            .akku_o_c_8(akku_o_c_8), .n46237(n46237), .n46211(n46211), 
            .n23757(n23757));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(43[10:18])
    \sram64kx8("sram64kx8.dat")(1,13)  RAM (.data({data}), .address({address}), 
            .data_7__N_89({data_7__N_89}), .akku_o_c_4(akku_o_c_4), .n46211(n46211), 
            .data_7__N_102(data_7__N_102), .n46237(n46237), .n23757(n23757), 
            .akku_o_c_0(akku_o_c_0), .akku_o_c_7(akku_o_c_7), .akku_o_c_6(akku_o_c_6), 
            .akku_o_c_5(akku_o_c_5), .akku_o_c_3(akku_o_c_3), .akku_o_c_2(akku_o_c_2), 
            .akku_o_c_1(akku_o_c_1), .reset_c(reset_c), .clk_c(clk_c), 
            .\states[0] (states[0]), .\states[1] (states[1]));   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(44[10:19])
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module CPU8BIT2
//

module CPU8BIT2 (states, clk_c, akku_o_c_0, address, data, GND_net, 
            akku_o_c_4, akku_o_c_1, akku_o_c_2, akku_o_c_3, \states[1] , 
            akku_o_c_7, data_7__N_89, data_7__N_102, akku_o_c_5, akku_o_c_6, 
            VCC_net, akku_o_c_8, n46237, n46211, n23757);
    output [2:0]states;
    input clk_c;
    output akku_o_c_0;
    output [5:0]address;
    input [7:0]data;
    input GND_net;
    output akku_o_c_4;
    output akku_o_c_1;
    output akku_o_c_2;
    output akku_o_c_3;
    output \states[1] ;
    output akku_o_c_7;
    input [7:0]data_7__N_89;
    input data_7__N_102;
    output akku_o_c_5;
    output akku_o_c_6;
    input VCC_net;
    output akku_o_c_8;
    output n46237;
    output n46211;
    output n23757;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(8[13:16])
    wire [8:0]n3;
    
    wire n45866;
    wire [4:0]n427;
    
    wire n45858, n46244;
    wire [2:0]states_2__N_76;
    
    wire n45850, n45848, n45856;
    wire [4:0]n640;
    
    wire n45843;
    wire [4:0]oprand;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(20[15:21])
    wire [9:0]n16;
    
    wire n46125, n43, n46870, n78, n46860, n45478;
    wire [5:0]adress_5__N_3;
    
    wire clk_c_enable_26, clk_c_enable_22;
    wire [8:0]n3555;
    
    wire n22545, n22535;
    wire [2:0]states_c;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(22[15:21])
    
    wire n22546;
    wire [5:0]pc;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(19[15:17])
    wire [5:0]pc_5__N_35;
    
    wire n22547, n22537, n22548, n46882, n7, n46121, n46136, n46060, 
        n45904, n46196, n38153, n22541, n22531, n22542, n46067, 
        n37, n46035, n46875, n46165, n45730, n45742, n45728, n45735, 
        n23094, n46850, n46307, n46068, n45978, n22543, n22533, 
        n22544, n41360, n22539, n22529, n22540, n40427;
    wire [5:0]n1012;
    wire [5:0]n1025;
    
    wire n46126;
    wire [8:0]n462;
    wire [8:0]n475;
    
    wire n44187, n44179;
    wire [8:0]n146;
    
    wire n55;
    wire [5:0]n2590;
    wire [8:0]n895;
    
    wire n43563, n46845, n182, n46028, n46029, n181, n211, n44171, 
        n44177, n45951, n44181, n46230;
    wire [5:0]n2577;
    
    wire n45749, n46058, n46037, n212, n46876, n6, n46878, n11, 
        n46266, n46108;
    wire [5:0]n1816;
    wire [8:0]n685;
    
    wire n89;
    wire [8:0]n720;
    
    wire n45787, n46017, n32, n43491, n43_adj_299, n46233, n46179, 
        n46064;
    wire [8:0]n218;
    
    wire n46090, n45976, n23881, n46155, n46057, n45844, n244, 
        n241, n243, n245, n45462, n583, n45865, n15, n46047, 
        n6_adj_300, n46309, n46310, n46370, n46844, n23, n43489, 
        n31, n23007, n46039, n46030, n169, n161, n191, n46880, 
        n37_adj_301, n45863, n22446, n45861, n45846, n40941, n43686, 
        n46143, n46852, n41054, n40006, n46034, n130, n160, n46020, 
        n41291, n43732, n45819, n8, n40426, n45847, n161_adj_302, 
        n43598, n43481, n51, n45724, n43706, n45727, n45725, n45474, 
        n46098, n22635, n45849, n46002, n46207, n46235, n22715, 
        n45786, n41378, n43532, n46857, n46858, n46859;
    wire [8:0]n112;
    
    wire n45390, n59, n45, n46085, n46056, n45987, n46027, n6324, 
        n45994, n46041, n46040;
    wire [8:0]n755;
    
    wire n45264;
    wire [5:0]n1543;
    wire [8:0]n615;
    
    wire n89_adj_303, n45794, n110, n106, n41356, n4, n45788, 
        n43595, n43479, n39, n40849, n41242, n45852, n45567, n46280, 
        n46281;
    wire [5:0]n2098;
    
    wire n46282;
    wire [5:0]n1324;
    
    wire n6_adj_304, n40788, n215, n117, n5, n117_adj_305, n10, 
        n43655, n38250, n46303, n46304, n46305, n118_adj_306, n46191, 
        n118_adj_307, n46163, n43668, n46264, n44022, n46006, n44765, 
        n44162, n46137, n45461;
    wire [8:0]n17;
    
    wire n45463, n46268, n87, n8_adj_310, n46225, n46229, n110_adj_311, 
        n106_adj_312, n41396, n31047, n29, n36, n39_adj_313, n2, 
        n40425, n46212, n46147, n45771, n45747, n46213, n87_adj_314, 
        n87_adj_315, n23565, n86, n43349;
    wire [8:0]n396;
    
    wire n45917, n15_adj_316, n45859, n4_adj_317, n46036, n45979, 
        mult_5u_5u_0_pp_2_6, n45968, n45596, n46214;
    wire [5:0]n2203;
    
    wire n43670, n45750, n40424;
    wire [5:0]n999;
    
    wire n14;
    wire [8:0]akku_o_8__N_50;
    
    wire n46854, n3622, n37_adj_318, n46019, n46168, n46240;
    wire [4:0]n1;
    
    wire n45853, n46300, n46301, n122, n40423, n46189, n46205, 
        n45851;
    wire [8:0]n790;
    
    wire n9081, n46270, mult_5u_5u_0_pp_2_5, mult_5u_5u_0_pp_2_4, mult_5u_5u_0_pp_1_2, 
        mult_5u_5u_0_cin_lr_2, co_mult_5u_5u_0_0_1, mult_5u_5u_0_pp_0_2, 
        co_mult_5u_5u_0_0_2, s_mult_5u_5u_0_0_4, mult_5u_5u_0_pp_0_4, 
        mult_5u_5u_0_pp_0_3, mult_5u_5u_0_pp_1_4, mult_5u_5u_0_pp_1_3, 
        co_mult_5u_5u_0_0_3, s_mult_5u_5u_0_0_5, s_mult_5u_5u_0_0_6, mult_5u_5u_0_pp_0_6, 
        mult_5u_5u_0_pp_0_5, mult_5u_5u_0_pp_1_6, mult_5u_5u_0_pp_1_5, 
        s_mult_5u_5u_0_0_7, s_mult_5u_5u_0_0_8, mult_5u_5u_0_pp_1_8, mult_5u_5u_0_pp_1_7, 
        co_t_mult_5u_5u_0_1_1, co_t_mult_5u_5u_0_1_2, mult_5u_5u_0_pp_2_7, 
        mult_5u_5u_0_pp_2_8, mult_5u_5u_0_cin_lr_0, mco, mco_1, mco_2, 
        mco_3, n46861, n46156, n46123, n43558, n43554, n83, n46049, 
        n46022, n22192;
    wire [2:0]n3668;
    
    wire n43750, n23490;
    wire [8:0]akku_o_8__N_67;
    
    wire n46276, n213, n46271, n40744, n40539, n22716, n46004;
    wire [8:0]n231;
    wire [8:0]n261;
    
    wire n45872;
    wire [4:0]n541;
    wire [8:0]n330;
    
    wire n45570, n40538, n40537, n45991, n45722, n46138, n45757;
    wire [8:0]n825;
    
    wire n43557, n31_adj_319, n46145, n89_adj_320, n46066, n46045, 
        n40422, n40536, n46021, n217;
    wire [8:0]n545;
    
    wire n45823, n45790;
    wire [5:0]n1687;
    
    wire n40740, n23044, n45822, n21753, n45892, n38297, n6_adj_321, 
        n7_adj_322, n40534, n46038, n46050, n46005, n117_adj_323;
    wire [8:0]n18;
    
    wire n44028, n43834, n221, n44030, n224, n45970, n40533;
    wire [8:0]n201;
    
    wire n40532, n46061, n46042, n46062, n46010, n40530, n4_adj_325, 
        n12, n45931, n191_adj_326, n45946, n45927, n45961;
    wire [8:0]n20;
    
    wire n40529, n45953, n41038, n45945, n45954, n46000, n40528, 
        n43883, n8_adj_331, n45975, n45952, n45943, n22712, n45965, 
        n45944, n40526, n22673, n45922, n221_adj_333, n220;
    wire [8:0]n270;
    
    wire n46296, n46297, n46873, n40525, n223, n222_adj_334, n191_adj_335, 
        n40524, n45932, n45916, n45925, n46223, n40523, n43353, 
        n45937, n107, n22035, n73_adj_336, n43333, n30878, n108, 
        n45997, n30783, n46173, n40522, n46197, n40521, n46199, 
        n46198, n40520, n46200, n46175, n40519, n46202, n46201, 
        n30723, n44099, n44026;
    wire [8:0]n270_adj_514;
    
    wire n46181;
    wire [7:0]n4247;
    
    wire n40518;
    wire [5:0]n2616;
    wire [5:0]n2629;
    
    wire n40517, n40516, n46120, n102, n22585, n46104, n45942, 
        n22969, n46111, n46044, n43707, n45285, n45284, n45286, 
        n8_adj_338, n46209;
    wire [8:0]n860;
    
    wire n40515;
    wire [5:0]n2603;
    
    wire n40514, n40513, n43712, n45731, n46157, n45738, n40512, 
        n40511, n40510, n43673, n7_adj_339, n45743, n40509, n40508, 
        n46096, n46083, n46097, n46851, n37_adj_340, n45862, n45908, 
        n45915, n43592, n45751, n6_adj_341, n8_adj_342;
    wire [4:0]n449;
    
    wire n45845, n46009, n39_adj_343, n51_adj_344, n45836, n168;
    wire [8:0]n363;
    
    wire n45816;
    wire [5:0]n2345;
    wire [4:0]n866;
    
    wire n51_adj_345, n43720, n43729;
    wire [5:0]n2358;
    
    wire n45864;
    wire [5:0]n2371;
    
    wire n46177, n46129, n40507, n43581, n46016;
    wire [4:0]n910;
    wire [8:0]n429;
    
    wire n257;
    wire [8:0]n208;
    
    wire n107_adj_346, n45287, n46171, n46261, n45481, n45807, n45929, 
        n45940, n45924, n40781, n19, n45923, n45914, n46114, n45762, 
        n45754, n43709, n43710, n43695, n22894, n41385, n40421, 
        n45900, n46409, n45933, n6383, n46110;
    wire [5:0]n2332;
    
    wire n45758, n4_adj_347, n4_adj_348, n21933, n9938, n44713, 
        n45732, n45726;
    wire [5:0]n2734;
    
    wire n44699;
    wire [5:0]n1855;
    
    wire n2_adj_349, n6_adj_350, n4_adj_351, n46848, n43759, n45867;
    wire [5:0]n2476;
    
    wire n46316, n46315, n43941, n45782;
    wire [8:0]n650;
    
    wire n45784, n45489;
    wire [8:0]n21;
    
    wire n46406, n46071, n29_adj_353, n45694, n46249, n43564, n46318, 
        n117_adj_354, n46320, n46319, n46323, n46322, n40506, n43991, 
        n6_adj_355, n2662, n46128, n45_adj_356, n46074, n45902, 
        n40960;
    wire [8:0]n231_adj_515;
    
    wire n4_adj_357, n10022, n22855;
    wire [4:0]n293;
    
    wire n21951, n46215, n109, n43606, n46403, n46385, n46379, 
        n46329, n45869, n46088, n12_adj_358, n152, n6_adj_359, n46332, 
        n46331, n46075, n46048, n45854, n46335, n46334, n46338, 
        n46337, n46025, n46089, n46078, n130_adj_360, n46091, n46183, 
        n46341, n40505;
    wire [4:0]n22564;
    
    wire n45778, n46130, n45773, n46340, n46344, n40504, n45776, 
        n45898, n41358, n45875, n6_adj_361, n46053, n46343, n160_adj_362, 
        n46351, n46350, n46354, n46353, n46073, n46357, n46356, 
        n46079, n46093, n46360, n46359, n45874, n45921, n22874, 
        n23447;
    wire [5:0]n2072;
    
    wire n46363, n46362, n46065, n46160, n46366, n46365, n46369, 
        n46400, n46368;
    wire [5:0]n1829;
    
    wire n46847, n46051, n45885, n46372, n45829, n46371, n4_adj_363, 
        n46375, n46378, n46084, n46381, n45974, n45981, n45982, 
        n46380, n46853, n21411, n46384, n46383, n46387, n46386, 
        n45729, n46390, n9, n40420, n43902, n30789, n46389, n46248, 
        n31204;
    wire [8:0]n930;
    
    wire n45475, n2_adj_367, n108_adj_368, n46396, n253, n256, n46395, 
        n45896, n46122, n6_adj_369, n45779;
    wire [5:0]n1051;
    
    wire n4_adj_370, n46399, n46398, n7_adj_371, n8_adj_372, n41383, 
        n6_adj_373, n77, n46402, n46293, n46294;
    wire [5:0]n1582;
    
    wire n4_adj_374, n46405, n45877, n45920, n43689, n46404, n122_adj_375, 
        n46288;
    wire [4:0]n405;
    
    wire n46408, n40419, n46287, n46407, n6_adj_376, n45909, n43766, 
        n43765, n45824, n6_adj_377, n22740, n6_adj_378, n9966, n21939, 
        n45753, n46086, n45842, n9959, n21937, n4_adj_379, n4_adj_380;
    wire [8:0]n580;
    wire [5:0]n1429;
    
    wire n45796, n45547, n43769, n11_adj_381, n9_adj_382, n22902, 
        n45870, n43768, n41077, n42171, n44079, n46087, n46059, 
        n41411, n45880, n22900, n41374, n6_adj_383, n41402, n4_adj_384, 
        n45918, n43675, n46055, n43547, n45871, n6734, n9_adj_385, 
        n45752, n4_adj_386, n45723, n45765, n45760, n45791, n40503, 
        n46069, n11_adj_388, n45663, n45912, n46397, n46052;
    wire [5:0]n1947;
    
    wire n45764, n23877, n45770, n45761, n46092, n46031, n23650, 
        n46082;
    wire [4:0]n4201;
    
    wire n45881;
    wire [5:0]n4217;
    
    wire n45883, n4_adj_389, n40857, n45876;
    wire [5:0]n2046;
    
    wire n40502, n2_adj_390, n46095, n45947;
    wire [5:0]n1842;
    
    wire n45763;
    wire [5:0]n2319;
    
    wire n40501, n7_adj_392, n45766, n40913, n45789, n45633, n4_adj_393, 
        n45899;
    wire [5:0]n2059;
    
    wire n8965, n45910, n45583, n46101, n45886, n45840, n45568, 
        n8_adj_394;
    wire [2:0]n4382;
    
    wire n45884, n45818, n45820, n45887, n45888;
    wire [5:0]n1403;
    
    wire n40970, n46100, n45626, n22924, n12_adj_395, n45566, n45878, 
        n23051, n46867, n45879, n38301, n45571, n46124, n45828, 
        n23030, n4_adj_396, n124, n46099, n40500, n45756, n45740, 
        n30, n43701, n7_adj_397, n45636, n45759, n6_adj_398, n23553, 
        n45733, n21510, n46243, n3611, n6_adj_399, n46033, n23541, 
        n45939, n45919, n45913, n45585, n8_adj_400, n23445, n43683, 
        n45769, n8_adj_401, n6_adj_402, n45800, n4_adj_403;
    wire [5:0]n4233;
    
    wire n22463;
    wire [5:0]n1156;
    
    wire n46043, n45806;
    wire [5:0]n1169;
    
    wire n46115, n30175, n46103;
    wire [3:0]n4330;
    
    wire n6_adj_404, n6574, n45873, n45985, n220_adj_405, n45966, 
        n45941, n45346, n7_adj_406, n45768, n6_adj_407, n22852, 
        n6_adj_408, n46102, n46118, n46077, n45936, n45901, n46081;
    wire [5:0]n1285;
    wire [5:0]n1416;
    
    wire n45868, n45855, n8_adj_409, n46003, n45620, n45827;
    wire [7:0]n4257;
    
    wire n40499, n45804, n46106, n6_adj_410, n46109, n23063, n21696, 
        n40498, n23806, n40497, n45830, n45734, n22479, n45627, 
        n6_adj_411, n40779, n21707, n5_adj_413, n40496, n23019, 
        n46866, n40495, n46146, n40494, n40493, n40492, clk_c_enable_20, 
        n45903, n46023, n190, n46112, n40830, n6_adj_414, n45894, 
        n46076, n45632, n46107, n67, n45889, n45634, n45890, n45891;
    wire [4:0]n4400;
    
    wire n41244, n5_adj_415, n43785, n6_adj_416, n45652, n45635, 
        n4_adj_417, n45905, n46869, n45906, n4_adj_418, n6_adj_419, 
        n8_adj_420, n43714, n22867, n7_adj_421, n41286, n45774, 
        n6_adj_422, n8_adj_423, n7_adj_424;
    wire [8:0]n270_adj_516;
    
    wire n45348, n46113, n45653, n45661, n255, n251, n254, n250, 
        n45662, n251_adj_429, n45956, n254_adj_430, n45950, n45351, 
        n45352, n46054, n46046, n21418, n6_adj_431, n21482, n23515, 
        n45928, n6_adj_432, n46116, n46117, n45907, n8_adj_433, 
        n22978, n45350, n45930, n45736, n46012, n45895, n41108, 
        n45821, n8_adj_434, n45860, n45973, n221_adj_435, n45972, 
        n45775, n23779, n45792, n45926, n45911, n5_adj_436;
    wire [4:0]n754;
    
    wire n122_adj_437, n15_adj_438, n13, n14_adj_439, n4_adj_440, 
        n46132, n23081, n45834, n21624, n7658, n43762, n45691, 
        n93, n45841, n41371, n21583, n6_adj_441, n46127, n46849, 
        n40491, n45777, n40490;
    wire [4:0]n4445;
    
    wire n23068, n45619, n40489, n45781, n8_adj_442, n820, n43753, 
        n7_adj_443, n45572, n45546, n5_adj_444, n40487, n4_adj_446, 
        n45999, n45983, n45998, n45969, n21395, n40486, n45988, 
        n45882, n46170, n46204, n40485, n8_adj_451, n46008, n45995, 
        n7_adj_452, n254_adj_453, n46382, n251_adj_454, n8_adj_455, 
        n43341, n45795, n45989, n250_adj_456, n46589, n248, n40484;
    wire [5:0]n2085;
    
    wire n40483, n40482, n12_adj_457, n30876, n246_adj_458, n242_adj_459, 
        n45935, n40417, n45949, n5_adj_460, n40481, n250_adj_461, 
        n6_adj_462, n40416;
    wire [8:0]n22;
    
    wire n40480, n46018, n45803, n40479, n23079, n30979, n40415, 
        n45971, n8_adj_464, n8_adj_465, n45799, n23659, n46133;
    wire [5:0]n1298;
    
    wire n45812, n41282, n45809, n6_adj_466, n43738, n46014, n45797, 
        n21590, n45832, n46151, n45802, n43678, n4_adj_467;
    wire [8:0]n510;
    
    wire n46144, n22998, n40801, n7458, n7_adj_468, n45801, n22887, 
        n7_adj_469, n43741, n6_adj_470, n45805, n7_adj_471, n8_adj_472;
    wire [4:0]n776;
    
    wire n41143, n40708, n30785, n45814, n40478, n46150, n46339, 
        n41354, n45785, n40477, n45957, n45958, n45825, n43727, 
        n40476, n45374;
    wire [5:0]n1038;
    
    wire n41388, n40475, n103, n46376, n40474, n40473, n45783;
    wire [5:0]n2293;
    
    wire n40413, n45964, n43679, n8_adj_476, n22896, n45793, n40472, 
        n46026, n45831, n40471, n40470, n46015, n8_adj_477, n45948, 
        n46164, n46364, n46166, n46167, n9_adj_478, n46790;
    wire [5:0]n2216;
    
    wire n46159, n43708, n45938, n23471, n40412, n21806, n21805;
    wire [5:0]n2489;
    
    wire n40411, n45992, n45963, n40410, n23070, n9_adj_484, n114, 
        n40469, n21777, n45741, n6_adj_485, n21776, n45833, n8_adj_486, 
        n9_adj_487, n40468, n45808, n41124, n46188;
    wire [3:0]n12888;
    
    wire n45780, n4_adj_488, n45491, n44729, n40467;
    wire [5:0]n1569;
    
    wire n43681, n4_adj_489, n40466, n40465, n45548, n8_adj_490;
    wire [5:0]n1311;
    
    wire n40464, n6_adj_491, n40463, n45986, n45960, n43647, n45739, 
        n45962, n13_adj_492, n159, n10_adj_493, n7_adj_494, n278_adj_495, 
        n40462, n15_adj_496, n45980, n40461, n40766, n4_adj_497, 
        n109_adj_498, n46345, n46324, n46330, n40460, n40459, n4_adj_499, 
        n46013, n45817, n45815, n41285, n40458, n43400, n46342, 
        n4_adj_500, n46001, n46206, n46210, n40457, n46336, n31179, 
        n46195, n40456, n40409, n46388, n45721, n21872, n40455, 
        n45955, n40454;
    wire [5:0]n1556;
    
    wire n46193, n45404, n40453, n40452, n31_adj_501, n46864, n45745, 
        n7_adj_502, n107_adj_503, n106_adj_504, n15_adj_505, n14_adj_506, 
        n30180, n46186, n30168, n40408, n46863, n45490, n40407, 
        n46257, n46258, n40451, n40450, n40449, n5_adj_507, n46245, 
        n46367, n46250, n46256, n40448, n12_adj_508, n46007, n45996, 
        n40447;
    wire [5:0]n1530;
    
    wire n40446, n38213, n6_adj_509, n45835, n40406, n45977, n40445, 
        n40444, n40405, n45248, n40443, n40442, n45984, n46277, 
        n122_adj_510, n46247, n45839, n40441, n45247, n45480, n66, 
        n40440, n45990, n122_adj_511, n117_adj_512, n40439, n40438, 
        n40437, n45838, n45810, n40436, n40435, n45479, n22207, 
        n46358, n40434, n22209, n22210, n4_adj_513, n40433, n40432, 
        n40431, n40430, n40429, n40428;
    
    LUT4 i2654_3_lut_rep_737_4_lut_4_lut_4_lut (.A(n3[3]), .B(n45866), .C(n3[2]), 
         .D(n427[1]), .Z(n45858)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (B (D)+!B (C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2654_3_lut_rep_737_4_lut_4_lut_4_lut.init = 16'hf710;
    FD1S3IX states__i0 (.D(states_2__N_76[0]), .CK(clk_c), .CD(n46244), 
            .Q(states[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam states__i0.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_722_4_lut (.A(n45850), .B(n45848), .C(n45856), .D(n640[1]), 
         .Z(n45843)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_rep_722_4_lut.init = 16'h718e;
    LUT4 i15268_2_lut_rep_1004_3_lut_3_lut_4_lut (.A(oprand[0]), .B(akku_o_c_0), 
         .C(n16[8]), .D(n16[7]), .Z(n46125)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam i15268_2_lut_rep_1004_3_lut_3_lut_4_lut.init = 16'h1e10;
    LUT4 i38124_2_lut_rep_1002_4_lut_else_3_lut (.A(n43), .B(n46870), .C(oprand[1]), 
         .D(n78), .Z(n46860)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i38124_2_lut_rep_1002_4_lut_else_3_lut.init = 16'hfffd;
    LUT4 oprand_3__bdd_4_lut_3_lut (.A(oprand[0]), .B(oprand[4]), .C(oprand[2]), 
         .Z(n45478)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam oprand_3__bdd_4_lut_3_lut.init = 16'h8080;
    FD1S3AX adreg_i0 (.D(adress_5__N_3[0]), .CK(clk_c), .Q(address[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam adreg_i0.GSR = "ENABLED";
    FD1P3AX oprand_i0_i0 (.D(data[0]), .SP(clk_c_enable_26), .CK(clk_c), 
            .Q(oprand[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam oprand_i0_i0.GSR = "ENABLED";
    FD1P3AX akku_i0_i1 (.D(n3555[0]), .SP(clk_c_enable_22), .CK(clk_c), 
            .Q(akku_o_c_0)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam akku_i0_i1.GSR = "ENABLED";
    PFUMX i15819 (.BLUT(n22545), .ALUT(n22535), .C0(states_c[2]), .Z(n22546));
    FD1P3AX pc_i0_i5 (.D(pc_5__N_35[5]), .SP(clk_c_enable_26), .CK(clk_c), 
            .Q(pc[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam pc_i0_i5.GSR = "ENABLED";
    PFUMX i15821 (.BLUT(n22547), .ALUT(n22537), .C0(states_c[2]), .Z(n22548));
    LUT4 i15282_2_lut_rep_1000_3_lut_4_lut (.A(n46882), .B(akku_o_c_0), 
         .C(n7), .D(n16[8]), .Z(n46121)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i15282_2_lut_rep_1000_3_lut_4_lut.init = 16'hfef0;
    LUT4 i31419_2_lut_3_lut_3_lut_4_lut (.A(n46136), .B(n46060), .C(n45904), 
         .D(n46196), .Z(n38153)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(C (D)))) */ ;
    defparam i31419_2_lut_3_lut_3_lut_4_lut.init = 16'h7000;
    PFUMX i15815 (.BLUT(n22541), .ALUT(n22531), .C0(states_c[2]), .Z(n22542));
    LUT4 i1_2_lut_rep_914_3_lut_4_lut (.A(n46067), .B(n37), .C(n46196), 
         .D(n46136), .Z(n46035)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_914_3_lut_4_lut.init = 16'h2000;
    LUT4 rem_59_i85_3_lut_rep_1044_4_lut_4_lut_4_lut (.A(oprand[2]), .B(n46875), 
         .C(oprand[1]), .D(oprand[4]), .Z(n46165)) /* synthesis lut_function=(A (C+!(D))+!A !((C+!(D))+!B)) */ ;
    defparam rem_59_i85_3_lut_rep_1044_4_lut_4_lut_4_lut.init = 16'ha4aa;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n45730), .B(n45742), .C(n45728), .D(n45735), 
         .Z(n23094)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hccc9;
    PFUMX i38446 (.BLUT(n46850), .ALUT(n46307), .C0(n46068), .Z(n45978));
    PFUMX i15817 (.BLUT(n22543), .ALUT(n22533), .C0(states_c[2]), .Z(n22544));
    LUT4 i1_2_lut_3_lut_4_lut (.A(n45850), .B(n45848), .C(n45856), .D(n640[1]), 
         .Z(n41360)) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hdb24;
    PFUMX i15813 (.BLUT(n22539), .ALUT(n22529), .C0(states_c[2]), .Z(n22540));
    CCU2D add_279_7 (.A0(n1012[4]), .B0(n1012[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40427), 
          .S0(n1025[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_279_7.INIT0 = 16'h5999;
    defparam add_279_7.INIT1 = 16'h0000;
    defparam add_279_7.INJECT1_0 = "NO";
    defparam add_279_7.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_1005_4_lut_3_lut_4_lut (.A(oprand[0]), .B(akku_o_c_0), 
         .C(n16[8]), .D(n16[7]), .Z(n46126)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i2_3_lut_rep_1005_4_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 mux_111_i4_3_lut_4_lut (.A(n46136), .B(n46060), .C(n46196), .D(n462[3]), 
         .Z(n475[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam mux_111_i4_3_lut_4_lut.init = 16'hf808;
    PFUMX i85 (.BLUT(n44187), .ALUT(n44179), .C0(n146[1]), .Z(n55));
    LUT4 mux_202_i5_3_lut_rep_1159 (.A(n2590[5]), .B(n895[4]), .C(n43563), 
         .Z(n46845)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_202_i5_3_lut_rep_1159.init = 16'h5c5c;
    LUT4 div_28_i147_3_lut_4_lut (.A(n182), .B(n46028), .C(n46029), .D(n181), 
         .Z(n211)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_i147_3_lut_4_lut.init = 16'hfe01;
    PFUMX i84 (.BLUT(n44171), .ALUT(n44177), .C0(n45951), .Z(n44181));
    LUT4 i1_2_lut_rep_1109_3_lut_4_lut (.A(oprand[1]), .B(n46882), .C(oprand[3]), 
         .D(oprand[2]), .Z(n46230)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_1109_3_lut_4_lut.init = 16'hfffe;
    LUT4 mux_202_i6_3_lut_rep_628 (.A(n2577[5]), .B(n895[5]), .C(n43563), 
         .Z(n45749)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_202_i6_3_lut_rep_628.init = 16'h5c5c;
    LUT4 div_28_i148_3_lut_4_lut_4_lut (.A(n46058), .B(n182), .C(n46029), 
         .D(n46037), .Z(n212)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B)) */ ;
    defparam div_28_i148_3_lut_4_lut_4_lut.init = 16'hccc6;
    LUT4 i32851_2_lut_3_lut (.A(oprand[1]), .B(n46882), .C(n46876), .Z(n6)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i32851_2_lut_3_lut.init = 16'hfefe;
    LUT4 i15147_2_lut_rep_987_3_lut_4_lut (.A(n46878), .B(n46882), .C(n11), 
         .D(n46266), .Z(n46108)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i15147_2_lut_rep_987_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i15758_2_lut_rep_666_4_lut (.A(n1816[5]), .B(n685[4]), .C(n89), 
         .D(n720[5]), .Z(n45787)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A (B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i15758_2_lut_rep_666_4_lut.init = 16'hff5c;
    LUT4 i38128_2_lut_rep_896_2_lut_3_lut_4_lut (.A(n46136), .B(n46060), 
         .C(n475[8]), .D(n46196), .Z(n46017)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C))+!A (C))) */ ;
    defparam i38128_2_lut_rep_896_2_lut_3_lut_4_lut.init = 16'h070f;
    PFUMX i55 (.BLUT(n32), .ALUT(n43491), .C0(akku_o_c_0), .Z(n43_adj_299));
    LUT4 i33082_2_lut_rep_1112_3_lut (.A(n46878), .B(n46882), .C(oprand[2]), 
         .Z(n46233)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i33082_2_lut_rep_1112_3_lut.init = 16'he0e0;
    LUT4 i1_2_lut_rep_855_4_lut_4_lut (.A(n46179), .B(n46064), .C(n218[5]), 
         .D(n46090), .Z(n45976)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(D))) */ ;
    defparam i1_2_lut_rep_855_4_lut_4_lut.init = 16'h7d28;
    LUT4 i32003_2_lut_rep_907_3_lut_4_lut_4_lut (.A(n46058), .B(n23881), 
         .C(n46155), .D(n46057), .Z(n46028)) /* synthesis lut_function=(!(A (B ((D)+!C)))) */ ;
    defparam i32003_2_lut_rep_907_3_lut_4_lut_4_lut.init = 16'h77f7;
    LUT4 i3085_3_lut_rep_723_4_lut (.A(n45850), .B(n45848), .C(n45856), 
         .D(n640[1]), .Z(n45844)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B ((D)+!C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3085_3_lut_rep_723_4_lut.init = 16'hdf04;
    LUT4 n264_bdd_4_lut (.A(n244), .B(n241), .C(n243), .D(n245), .Z(n45462)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n264_bdd_4_lut.init = 16'hfffe;
    LUT4 mux_86_i4_3_lut_rep_727 (.A(n583), .B(n45865), .C(n15), .Z(n45848)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_86_i4_3_lut_rep_727.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut (.A(n23881), .B(n46047), .C(n46029), .D(n212), 
         .Z(n6_adj_300)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_4_lut.init = 16'hff56;
    LUT4 n46309_bdd_4_lut (.A(n46309), .B(n46310), .C(akku_o_c_4), .D(n46370), 
         .Z(n46844)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n46309_bdd_4_lut.init = 16'hca00;
    PFUMX i54 (.BLUT(n23), .ALUT(n43489), .C0(oprand[0]), .Z(n31));
    LUT4 i1_2_lut_3_lut_4_lut_adj_74 (.A(n46136), .B(n46060), .C(n475[8]), 
         .D(n46196), .Z(n23007)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_74.init = 16'h78f0;
    LUT4 div_39_i133_3_lut_4_lut (.A(n46039), .B(n46030), .C(n169), .D(n161), 
         .Z(n191)) /* synthesis lut_function=(A (B (D)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_i133_3_lut_4_lut.init = 16'hf807;
    LUT4 mux_22_i8_3_lut_rep_1015_4_lut (.A(oprand[0]), .B(n46880), .C(n16[8]), 
         .D(n16[7]), .Z(n46136)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_22_i8_3_lut_rep_1015_4_lut.init = 16'hfe10;
    LUT4 i3243_2_lut_4_lut (.A(n45850), .B(n45856), .C(n37_adj_301), .D(n45863), 
         .Z(n22446)) /* synthesis lut_function=(A (B+(C+!(D)))+!A !(B (C (D))+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i3243_2_lut_4_lut.init = 16'hacff;
    LUT4 i3230_2_lut_rep_725_4_lut (.A(n45850), .B(n45856), .C(n37_adj_301), 
         .D(n45861), .Z(n45846)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i3230_2_lut_rep_725_4_lut.init = 16'h53ac;
    LUT4 i1_2_lut_rep_729 (.A(n40941), .B(n43686), .Z(n45850)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_rep_729.init = 16'h6666;
    LUT4 i1_2_lut_2_lut_3_lut (.A(n46143), .B(n46852), .C(n46155), .Z(n41054)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;
    defparam i1_2_lut_2_lut_3_lut.init = 16'h6969;
    LUT4 i33272_2_lut_3_lut (.A(akku_o_c_1), .B(akku_o_c_0), .C(akku_o_c_2), 
         .Z(n40006)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i33272_2_lut_3_lut.init = 16'h8080;
    LUT4 i24525_3_lut_2_lut_3_lut_4_lut (.A(n46068), .B(n46034), .C(n130), 
         .D(n46850), .Z(n160)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i24525_3_lut_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i32011_2_lut_rep_899_3_lut_4_lut_4_lut (.A(n46058), .B(n182), .C(n46047), 
         .D(n23881), .Z(n46020)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;
    defparam i32011_2_lut_rep_899_3_lut_4_lut_4_lut.init = 16'hfdff;
    LUT4 i2_3_lut_rep_698_4_lut (.A(n40941), .B(n43686), .C(n41291), .D(n43732), 
         .Z(n45819)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i2_3_lut_rep_698_4_lut.init = 16'h6996;
    LUT4 i33054_2_lut_3_lut_4_lut (.A(akku_o_c_1), .B(n46880), .C(akku_o_c_3), 
         .D(akku_o_c_2), .Z(n8)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i33054_2_lut_3_lut_4_lut.init = 16'hfff8;
    CCU2D add_279_5 (.A0(n1012[2]), .B0(n1012[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1012[3]), .B1(n1012[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40426), .COUT(n40427), .S0(n1025[3]), .S1(n1025[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_279_5.INIT0 = 16'h5999;
    defparam add_279_5.INIT1 = 16'h5666;
    defparam add_279_5.INJECT1_0 = "NO";
    defparam add_279_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_1145 (.A(n46880), .B(akku_o_c_1), .Z(n46266)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1145.init = 16'heeee;
    LUT4 i3078_4_lut_3_lut_rep_726_4_lut (.A(n40941), .B(n43686), .C(n45856), 
         .D(n45848), .Z(n45847)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C+!(D))))) */ ;
    defparam i3078_4_lut_3_lut_rep_726_4_lut.init = 16'h6f06;
    LUT4 div_53_i112_3_lut_4_lut_3_lut_4_lut (.A(n46068), .B(n46034), .C(n130), 
         .D(n46850), .Z(n161_adj_302)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_i112_3_lut_4_lut_3_lut_4_lut.init = 16'h7780;
    PFUMX i63 (.BLUT(n43598), .ALUT(n43481), .C0(n46880), .Z(n51));
    LUT4 n937_bdd_4_lut (.A(n45724), .B(n43706), .C(n45727), .D(n45725), 
         .Z(n45474)) /* synthesis lut_function=(A (B+(C+(D)))+!A ((C+!(D))+!B)) */ ;
    defparam n937_bdd_4_lut.init = 16'hfbfd;
    LUT4 i2_3_lut_4_lut (.A(n46136), .B(n46067), .C(n46098), .D(n46090), 
         .Z(n22635)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_93_i5_3_lut_rep_728_4_lut (.A(n40941), .B(n43686), .C(n37_adj_301), 
         .D(n45856), .Z(n45849)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_93_i5_3_lut_rep_728_4_lut.init = 16'h6f60;
    LUT4 i24524_2_lut_rep_881_3_lut_4_lut (.A(n46068), .B(n46034), .C(n130), 
         .D(n46850), .Z(n46002)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i24524_2_lut_rep_881_3_lut_4_lut.init = 16'hf8f0;
    LUT4 equal_1847_i7_2_lut_rep_1086_3_lut_4_lut (.A(n46880), .B(akku_o_c_1), 
         .C(n46882), .D(n46878), .Z(n46207)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam equal_1847_i7_2_lut_rep_1086_3_lut_4_lut.init = 16'hfffe;
    LUT4 i33575_2_lut_rep_1114_3_lut (.A(n46880), .B(akku_o_c_1), .C(akku_o_c_2), 
         .Z(n46235)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i33575_2_lut_rep_1114_3_lut.init = 16'he0e0;
    LUT4 i3_4_lut_4_lut (.A(n46058), .B(n182), .C(n181), .D(n23881), 
         .Z(n22715)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;
    defparam i3_4_lut_4_lut.init = 16'hfdff;
    LUT4 i15132_2_lut_rep_665_4_lut (.A(n1816[5]), .B(n685[4]), .C(n89), 
         .D(n720[5]), .Z(n45786)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B (D)+!B ((D)+!C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i15132_2_lut_rep_665_4_lut.init = 16'hffa3;
    LUT4 mux_22_i4_3_lut_rep_1034_4_lut (.A(n46882), .B(n46880), .C(n16[4]), 
         .D(n16[3]), .Z(n46155)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_22_i4_3_lut_rep_1034_4_lut.init = 16'hfe10;
    LUT4 i2_3_lut_4_lut_adj_75 (.A(n40941), .B(n43686), .C(n45856), .D(n45848), 
         .Z(n41378)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i2_3_lut_4_lut_adj_75.init = 16'h6996;
    LUT4 i2_3_lut_4_lut_3_lut (.A(akku_o_c_0), .B(akku_o_c_3), .C(akku_o_c_2), 
         .Z(n43532)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut_4_lut_3_lut.init = 16'h8080;
    PFUMX i38758 (.BLUT(n46857), .ALUT(n46858), .C0(akku_o_c_1), .Z(n46859));
    LUT4 mux_29_i4_3_lut_4_lut_4_lut (.A(n46155), .B(n46057), .C(n7), 
         .D(n22715), .Z(n112[3])) /* synthesis lut_function=(A ((C+(D))+!B)+!A !(C+!(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_29_i4_3_lut_4_lut_4_lut.init = 16'hafa2;
    FD1P3AX oprand_i0_i0_rep_1181 (.D(data[0]), .SP(clk_c_enable_26), .CK(clk_c), 
            .Q(n46882)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam oprand_i0_i0_rep_1181.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(n45390), .B(n59), .Z(n45)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i2213_2_lut_3_lut_4_lut_4_lut (.A(n46085), .B(n46056), .C(n45987), 
         .D(n46027), .Z(n6324)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2213_2_lut_3_lut_4_lut_4_lut.init = 16'h1000;
    LUT4 div_53_i113_3_lut_rep_873_4_lut_4_lut (.A(n46068), .B(n46034), 
         .C(n46850), .D(n130), .Z(n45994)) /* synthesis lut_function=(!(A (B (C+(D)))+!A !(B (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_i113_3_lut_rep_873_4_lut_4_lut.init = 16'h662a;
    LUT4 n758_bdd_3_lut_4_lut (.A(n46090), .B(n46041), .C(n46040), .D(n755[6]), 
         .Z(n45264)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(C+(D))) */ ;
    defparam n758_bdd_3_lut_4_lut.init = 16'h8887;
    LUT4 mux_146_i5_3_lut_rep_673 (.A(n1543[5]), .B(n615[4]), .C(n89_adj_303), 
         .Z(n45794)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_146_i5_3_lut_rep_673.init = 16'h5c5c;
    LUT4 i1_4_lut (.A(n110), .B(n106), .C(n41356), .D(n4), .Z(n43489)) /* synthesis lut_function=(!((B (C+!(D))+!B (C+(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_4_lut.init = 16'h0802;
    LUT4 i4609_2_lut_rep_667_4_lut (.A(n1816[5]), .B(n685[4]), .C(n89), 
         .D(n720[5]), .Z(n45788)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (D)+!B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i4609_2_lut_rep_667_4_lut.init = 16'h5c00;
    PFUMX i62 (.BLUT(n43595), .ALUT(n43479), .C0(n46882), .Z(n39));
    LUT4 mux_22_i5_3_lut_rep_1022_4_lut (.A(n46882), .B(n46880), .C(n16[5]), 
         .D(n16[4]), .Z(n46143)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_22_i5_3_lut_rep_1022_4_lut.init = 16'hfe10;
    LUT4 n41077_bdd_3_lut_4_lut (.A(n40849), .B(n41242), .C(n45852), .D(n45858), 
         .Z(n45567)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam n41077_bdd_3_lut_4_lut.init = 16'h23dc;
    PFUMX i38429 (.BLUT(n46280), .ALUT(n46281), .C0(n2098[3]), .Z(n46282));
    LUT4 i2_4_lut_4_lut (.A(n1324[3]), .B(n1324[5]), .C(n6_adj_304), .D(n1324[4]), 
         .Z(n40788)) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_4_lut_4_lut.init = 16'hdb24;
    LUT4 div_28_i151_3_lut_4_lut_4_lut_4_lut (.A(n46155), .B(n46057), .C(n22715), 
         .D(n41054), .Z(n215)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_i151_3_lut_4_lut_4_lut_4_lut.init = 16'hf301;
    LUT4 i3_4_lut (.A(n117), .B(n5), .C(n117_adj_305), .D(n10), .Z(n43655)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i31516_2_lut_3_lut_3_lut_4_lut (.A(n46090), .B(n46041), .C(n755[6]), 
         .D(n46040), .Z(n38250)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;
    defparam i31516_2_lut_3_lut_3_lut_4_lut.init = 16'h0070;
    PFUMX i38444 (.BLUT(n46303), .ALUT(n46304), .C0(akku_o_c_0), .Z(n46305));
    LUT4 i3_4_lut_adj_76 (.A(n118_adj_306), .B(n46191), .C(n118_adj_307), 
         .D(n46163), .Z(n43668)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i3_4_lut_adj_76.init = 16'hfffe;
    LUT4 i1_2_lut_rep_1143 (.A(n46878), .B(n46882), .Z(n46264)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_1143.init = 16'heeee;
    LUT4 i37135_2_lut_3_lut_4_lut (.A(n46090), .B(n46041), .C(n755[6]), 
         .D(n46040), .Z(n44022)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i37135_2_lut_3_lut_4_lut.init = 16'hfff8;
    LUT4 i1_2_lut_rep_885_4_lut (.A(n112[6]), .B(n112[4]), .C(n46207), 
         .D(n169), .Z(n46006)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_885_4_lut.init = 16'h35ca;
    LUT4 i38096_2_lut_rep_1016_3_lut_4_lut (.A(n46882), .B(n46880), .C(n44765), 
         .D(n44162), .Z(n46137)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i38096_2_lut_rep_1016_3_lut_4_lut.init = 16'hfffe;
    PFUMX i38298 (.BLUT(n45462), .ALUT(n45461), .C0(n17[1]), .Z(n45463));
    LUT4 i37117_2_lut_rep_1147 (.A(akku_o_c_3), .B(akku_o_c_2), .Z(n46268)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i37117_2_lut_rep_1147.init = 16'heeee;
    LUT4 rem_36_i63_3_lut_4_lut_3_lut (.A(akku_o_c_3), .B(akku_o_c_2), .C(akku_o_c_4), 
         .Z(n87)) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam rem_36_i63_3_lut_4_lut_3_lut.init = 16'h8a8a;
    LUT4 i6222_1_lut_3_lut_4_lut (.A(oprand[0]), .B(akku_o_c_0), .C(n16[4]), 
         .D(n16[3]), .Z(n8_adj_310)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B (C)))) */ ;
    defparam i6222_1_lut_3_lut_4_lut.init = 16'h01ef;
    LUT4 i24353_2_lut_rep_1104_3_lut_4_lut (.A(akku_o_c_3), .B(akku_o_c_2), 
         .C(akku_o_c_0), .D(akku_o_c_1), .Z(n46225)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i24353_2_lut_rep_1104_3_lut_4_lut.init = 16'hfeee;
    LUT4 i2_2_lut_rep_1108_3_lut_4_lut (.A(akku_o_c_3), .B(akku_o_c_2), 
         .C(akku_o_c_1), .D(n46880), .Z(n46229)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_2_lut_rep_1108_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_77 (.A(n110_adj_311), .B(n106_adj_312), .C(n41396), 
         .D(n31047), .Z(n43491)) /* synthesis lut_function=(!((B (C+!(D))+!B (C+(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_4_lut_adj_77.init = 16'h0802;
    PFUMX i62_adj_78 (.BLUT(n29), .ALUT(n36), .C0(n46882), .Z(n39_adj_313));
    LUT4 i5759_4_lut_4_lut (.A(n1324[2]), .B(n1324[5]), .C(n1324[1]), 
         .D(n2), .Z(n6_adj_304)) /* synthesis lut_function=(A ((C (D))+!B)+!A !(B+!(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5759_4_lut_4_lut.init = 16'hb332;
    CCU2D add_279_3 (.A0(n1012[0]), .B0(n1012[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1012[1]), .B1(n1012[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40425), .COUT(n40426), .S0(n1025[1]), .S1(n1025[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_279_3.INIT0 = 16'h5999;
    defparam add_279_3.INIT1 = 16'h5999;
    defparam add_279_3.INJECT1_0 = "NO";
    defparam add_279_3.INJECT1_1 = "NO";
    LUT4 i38163_2_lut_rep_1026_2_lut_3_lut_4_lut_4_lut (.A(akku_o_c_3), .B(akku_o_c_2), 
         .C(n46212), .D(akku_o_c_4), .Z(n46147)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C+(D)))+!A (B (C+!(D))+!B (C)))) */ ;
    defparam i38163_2_lut_rep_1026_2_lut_3_lut_4_lut_4_lut.init = 16'h0d03;
    LUT4 i5414_2_lut_rep_626_4_lut (.A(n2577[5]), .B(n895[5]), .C(n43563), 
         .D(n45771), .Z(n45747)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(B (D)+!B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i5414_2_lut_rep_626_4_lut.init = 16'ha35c;
    LUT4 i1_2_lut_rep_1092_3_lut (.A(akku_o_c_3), .B(akku_o_c_2), .C(akku_o_c_4), 
         .Z(n46213)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i1_2_lut_rep_1092_3_lut.init = 16'he0e0;
    LUT4 i3_4_lut_adj_79 (.A(n87_adj_314), .B(n87_adj_315), .C(n23565), 
         .D(n86), .Z(n43349)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i3_4_lut_adj_79.init = 16'hfffe;
    LUT4 mux_100_i6_3_lut_rep_738_4_lut (.A(n396[7]), .B(n45917), .C(n45863), 
         .D(n15_adj_316), .Z(n45859)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam mux_100_i6_3_lut_rep_738_4_lut.init = 16'hf080;
    LUT4 i2201_3_lut_rep_858_4_lut (.A(n4_adj_317), .B(n46036), .C(n45987), 
         .D(n46056), .Z(n45979)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !((D)+!C)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2201_3_lut_rep_858_4_lut.init = 16'h80f8;
    LUT4 i1983_1_lut (.A(address[0]), .Z(pc_5__N_35[0])) /* synthesis lut_function=(!(A)) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i1983_1_lut.init = 16'h5555;
    AND2 AND2_t2 (.A(akku_o_c_2), .B(oprand[4]), .Z(mult_5u_5u_0_pp_2_6)) /* synthesis syn_instantiated=1 */ ;   // mult_5u_5u.v(69[10:63])
    CCU2D add_279_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n46060), .B1(n46136), .C1(n46196), .D1(n462[3]), .COUT(n40425), 
          .S1(n1025[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_279_1.INIT0 = 16'hF000;
    defparam add_279_1.INIT1 = 16'h07f7;
    defparam add_279_1.INJECT1_0 = "NO";
    defparam add_279_1.INJECT1_1 = "NO";
    LUT4 i2208_3_lut_rep_847_4_lut_4_lut (.A(n46085), .B(n46056), .C(n45987), 
         .D(n46027), .Z(n45968)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B !(C+!(D))))) */ ;
    defparam i2208_3_lut_rep_847_4_lut_4_lut.init = 16'h10fb;
    LUT4 n398_bdd_4_lut_4_lut (.A(n396[7]), .B(n45917), .C(n45863), .D(n45849), 
         .Z(n45596)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A !(C (D))) */ ;
    defparam n398_bdd_4_lut_4_lut.init = 16'ha5d5;
    LUT4 i1_2_lut_rep_1093_3_lut (.A(akku_o_c_3), .B(akku_o_c_2), .C(akku_o_c_4), 
         .Z(n46214)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_1093_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_rep_629 (.A(n2203[5]), .B(n43670), .Z(n45750)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_rep_629.init = 16'h6666;
    CCU2D add_277_7 (.A0(n999[4]), .B0(n999[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40424), 
          .S0(n1012[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_277_7.INIT0 = 16'h5999;
    defparam add_277_7.INIT1 = 16'h0000;
    defparam add_277_7.INJECT1_0 = "NO";
    defparam add_277_7.INJECT1_1 = "NO";
    LUT4 i29_2_lut (.A(akku_o_c_3), .B(akku_o_c_4), .Z(n14)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    defparam i29_2_lut.init = 16'h6666;
    LUT4 i15808_4_lut (.A(akku_o_8__N_50[4]), .B(n45730), .C(n46854), 
         .D(n3622), .Z(n22535)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(73[13] 82[22])
    defparam i15808_4_lut.init = 16'hca0a;
    LUT4 mux_65_i7_3_lut_rep_898_4_lut (.A(n4_adj_317), .B(n46036), .C(n37_adj_318), 
         .D(n46056), .Z(n46019)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_65_i7_3_lut_rep_898_4_lut.init = 16'h8f80;
    LUT4 i33676_2_lut_rep_1047_3_lut_3_lut_4_lut (.A(akku_o_c_3), .B(akku_o_c_2), 
         .C(akku_o_c_4), .D(akku_o_c_1), .Z(n46168)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;
    defparam i33676_2_lut_rep_1047_3_lut_3_lut_4_lut.init = 16'h0fe0;
    LUT4 states_2__bdd_3_lut (.A(states_c[2]), .B(states[0]), .C(\states[1] ), 
         .Z(clk_c_enable_22)) /* synthesis lut_function=(!(A (B)+!A !(C))) */ ;
    defparam states_2__bdd_3_lut.init = 16'h7272;
    LUT4 i1_2_lut_rep_1119_3_lut (.A(akku_o_c_3), .B(akku_o_c_2), .C(akku_o_c_4), 
         .Z(n46240)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i1_2_lut_rep_1119_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_3_lut_4_lut_adj_80 (.A(n4_adj_317), .B(n46036), .C(n46056), 
         .D(n45987), .Z(n1[1])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_3_lut_4_lut_adj_80.init = 16'h7887;
    LUT4 i14914_3_lut_rep_732 (.A(n3[2]), .B(n41242), .C(n3[1]), .Z(n45853)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i14914_3_lut_rep_732.init = 16'h5151;
    PFUMX i38442 (.BLUT(n46300), .ALUT(n46301), .C0(akku_o_c_4), .Z(n122));
    CCU2D add_277_5 (.A0(n999[2]), .B0(n999[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n999[3]), .B1(n999[5]), .C1(GND_net), .D1(GND_net), .CIN(n40423), 
          .COUT(n40424), .S0(n1012[3]), .S1(n1012[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_277_5.INIT0 = 16'h5999;
    defparam add_277_5.INIT1 = 16'h5666;
    defparam add_277_5.INJECT1_0 = "NO";
    defparam add_277_5.INJECT1_1 = "NO";
    LUT4 i24313_2_lut_rep_1068_3_lut_4_lut (.A(akku_o_c_3), .B(akku_o_c_2), 
         .C(akku_o_c_1), .D(akku_o_c_4), .Z(n46189)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;
    defparam i24313_2_lut_rep_1068_3_lut_4_lut.init = 16'h70f0;
    LUT4 i2683_3_lut_rep_731_3_lut (.A(n3[2]), .B(n41242), .C(n3[1]), 
         .Z(n45852)) /* synthesis lut_function=(!(A (B+!(C))+!A !((C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2683_3_lut_rep_731_3_lut.init = 16'h7171;
    LUT4 i1_2_lut_3_lut (.A(akku_o_c_3), .B(akku_o_c_2), .C(akku_o_c_4), 
         .Z(n86)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h7070;
    LUT4 akku_o_c_2_bdd_3_lut_38408_rep_1084_4_lut_4_lut (.A(akku_o_c_3), 
         .B(akku_o_c_2), .C(akku_o_c_1), .D(akku_o_c_4), .Z(n46205)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B))) */ ;
    defparam akku_o_c_2_bdd_3_lut_38408_rep_1084_4_lut_4_lut.init = 16'h4ccc;
    LUT4 i14912_3_lut_rep_730_4_lut_4_lut (.A(n3[2]), .B(n41242), .C(n3[1]), 
         .D(n40849), .Z(n45851)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i14912_3_lut_rep_730_4_lut_4_lut.init = 16'h00fd;
    LUT4 i4970_2_lut_3_lut (.A(n2203[5]), .B(n43670), .C(n790[2]), .Z(n9081)) /* synthesis lut_function=(A (B (C))+!A !(B+!(C))) */ ;
    defparam i4970_2_lut_3_lut.init = 16'h9090;
    LUT4 i1_2_lut_rep_1149 (.A(akku_o_c_3), .B(akku_o_c_2), .C(akku_o_c_4), 
         .Z(n46270)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_1149.init = 16'h8080;
    AND2 AND2_t3 (.A(akku_o_c_1), .B(oprand[4]), .Z(mult_5u_5u_0_pp_2_5)) /* synthesis syn_instantiated=1 */ ;   // mult_5u_5u.v(67[10:63])
    AND2 AND2_t4 (.A(akku_o_c_0), .B(oprand[4]), .Z(mult_5u_5u_0_pp_2_4)) /* synthesis syn_instantiated=1 */ ;   // mult_5u_5u.v(65[10:63])
    AND2 AND2_t5 (.A(akku_o_c_0), .B(oprand[2]), .Z(mult_5u_5u_0_pp_1_2)) /* synthesis syn_instantiated=1 */ ;   // mult_5u_5u.v(63[10:63])
    AND2 AND2_t6 (.A(n46880), .B(n46882), .Z(n16[0])) /* synthesis syn_instantiated=1 */ ;   // mult_5u_5u.v(61[10:63])
    FADD2B mult_5u_5u_0_cin_lr_add_2 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_5u_5u_0_cin_lr_2)) /* synthesis syn_instantiated=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(35[23:37])
    FADD2B Cadd_mult_5u_5u_0_0_1 (.A0(GND_net), .A1(mult_5u_5u_0_pp_0_2), 
           .B0(GND_net), .B1(mult_5u_5u_0_pp_1_2), .CI(GND_net), .COUT(co_mult_5u_5u_0_0_1), 
           .S1(n16[2])) /* synthesis syn_instantiated=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(35[23:37])
    FADD2B mult_5u_5u_0_add_0_2 (.A0(mult_5u_5u_0_pp_0_3), .A1(mult_5u_5u_0_pp_0_4), 
           .B0(mult_5u_5u_0_pp_1_3), .B1(mult_5u_5u_0_pp_1_4), .CI(co_mult_5u_5u_0_0_1), 
           .COUT(co_mult_5u_5u_0_0_2), .S0(n16[3]), .S1(s_mult_5u_5u_0_0_4)) /* synthesis syn_instantiated=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(35[23:37])
    FADD2B mult_5u_5u_0_add_0_3 (.A0(mult_5u_5u_0_pp_0_5), .A1(mult_5u_5u_0_pp_0_6), 
           .B0(mult_5u_5u_0_pp_1_5), .B1(mult_5u_5u_0_pp_1_6), .CI(co_mult_5u_5u_0_0_2), 
           .COUT(co_mult_5u_5u_0_0_3), .S0(s_mult_5u_5u_0_0_5), .S1(s_mult_5u_5u_0_0_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(35[23:37])
    FADD2B mult_5u_5u_0_add_0_4 (.A0(GND_net), .A1(GND_net), .B0(mult_5u_5u_0_pp_1_7), 
           .B1(mult_5u_5u_0_pp_1_8), .CI(co_mult_5u_5u_0_0_3), .S0(s_mult_5u_5u_0_0_7), 
           .S1(s_mult_5u_5u_0_0_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(35[23:37])
    FADD2B Cadd_t_mult_5u_5u_0_1_1 (.A0(GND_net), .A1(s_mult_5u_5u_0_0_4), 
           .B0(GND_net), .B1(mult_5u_5u_0_pp_2_4), .CI(GND_net), .COUT(co_t_mult_5u_5u_0_1_1), 
           .S1(n16[4])) /* synthesis syn_instantiated=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(35[23:37])
    FADD2B t_mult_5u_5u_0_add_1_2 (.A0(s_mult_5u_5u_0_0_5), .A1(s_mult_5u_5u_0_0_6), 
           .B0(mult_5u_5u_0_pp_2_5), .B1(mult_5u_5u_0_pp_2_6), .CI(co_t_mult_5u_5u_0_1_1), 
           .COUT(co_t_mult_5u_5u_0_1_2), .S0(n16[5]), .S1(n16[6])) /* synthesis syn_instantiated=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(35[23:37])
    FADD2B t_mult_5u_5u_0_add_1_3 (.A0(s_mult_5u_5u_0_0_7), .A1(s_mult_5u_5u_0_0_8), 
           .B0(mult_5u_5u_0_pp_2_7), .B1(mult_5u_5u_0_pp_2_8), .CI(co_t_mult_5u_5u_0_1_2), 
           .S0(n16[7]), .S1(n16[8])) /* synthesis syn_instantiated=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(35[23:37])
    MULT2 mult_5u_5u_0_mult_0_0 (.A0(n46880), .A1(akku_o_c_1), .A2(akku_o_c_1), 
          .A3(akku_o_c_2), .B0(n46878), .B1(n46882), .B2(n46878), .B3(n46882), 
          .CI(mult_5u_5u_0_cin_lr_0), .CO(mco), .P0(n16[1]), .P1(mult_5u_5u_0_pp_0_2)) /* synthesis syn_instantiated=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(35[23:37])
    MULT2 mult_5u_5u_0_mult_0_1 (.A0(akku_o_c_2), .A1(akku_o_c_3), .A2(akku_o_c_3), 
          .A3(akku_o_c_4), .B0(oprand[1]), .B1(oprand[0]), .B2(oprand[1]), 
          .B3(oprand[0]), .CI(mco), .CO(mco_1), .P0(mult_5u_5u_0_pp_0_3), 
          .P1(mult_5u_5u_0_pp_0_4)) /* synthesis syn_instantiated=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(35[23:37])
    MULT2 mult_5u_5u_0_mult_0_2 (.A0(akku_o_c_4), .A1(GND_net), .A2(GND_net), 
          .A3(GND_net), .B0(oprand[1]), .B1(oprand[0]), .B2(oprand[1]), 
          .B3(oprand[0]), .CI(mco_1), .P0(mult_5u_5u_0_pp_0_5), .P1(mult_5u_5u_0_pp_0_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(35[23:37])
    MULT2 mult_5u_5u_0_mult_2_0 (.A0(akku_o_c_0), .A1(akku_o_c_1), .A2(akku_o_c_1), 
          .A3(akku_o_c_2), .B0(oprand[3]), .B1(oprand[2]), .B2(oprand[3]), 
          .B3(oprand[2]), .CI(mult_5u_5u_0_cin_lr_2), .CO(mco_2), .P0(mult_5u_5u_0_pp_1_3), 
          .P1(mult_5u_5u_0_pp_1_4)) /* synthesis syn_instantiated=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(35[23:37])
    MULT2 mult_5u_5u_0_mult_2_1 (.A0(akku_o_c_2), .A1(akku_o_c_3), .A2(akku_o_c_3), 
          .A3(akku_o_c_4), .B0(oprand[3]), .B1(oprand[2]), .B2(oprand[3]), 
          .B3(oprand[2]), .CI(mco_2), .CO(mco_3), .P0(mult_5u_5u_0_pp_1_5), 
          .P1(mult_5u_5u_0_pp_1_6)) /* synthesis syn_instantiated=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(35[23:37])
    MULT2 mult_5u_5u_0_mult_2_2 (.A0(akku_o_c_4), .A1(GND_net), .A2(GND_net), 
          .A3(GND_net), .B0(oprand[3]), .B1(oprand[2]), .B2(oprand[3]), 
          .B3(oprand[2]), .CI(mco_3), .P0(mult_5u_5u_0_pp_1_7), .P1(mult_5u_5u_0_pp_1_8)) /* synthesis syn_instantiated=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(35[23:37])
    AND2 AND2_t1 (.A(akku_o_c_3), .B(oprand[4]), .Z(mult_5u_5u_0_pp_2_7)) /* synthesis syn_instantiated=1 */ ;   // mult_5u_5u.v(71[10:63])
    AND2 AND2_t0 (.A(akku_o_c_4), .B(oprand[4]), .Z(mult_5u_5u_0_pp_2_8)) /* synthesis syn_instantiated=1 */ ;   // mult_5u_5u.v(73[10:63])
    FADD2B mult_5u_5u_0_cin_lr_add_0 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_5u_5u_0_cin_lr_0)) /* synthesis syn_instantiated=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(35[23:37])
    FD1P3AX pc_i0_i4 (.D(pc_5__N_35[4]), .SP(clk_c_enable_26), .CK(clk_c), 
            .Q(pc[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam pc_i0_i4.GSR = "ENABLED";
    PFUMX i38760 (.BLUT(n46860), .ALUT(n46861), .C0(n46156), .Z(n46123));
    FD1P3AX pc_i0_i3 (.D(pc_5__N_35[3]), .SP(clk_c_enable_26), .CK(clk_c), 
            .Q(pc[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam pc_i0_i3.GSR = "ENABLED";
    PFUMX i113 (.BLUT(n43558), .ALUT(n43554), .C0(n46876), .Z(n83));
    FD1P3AX pc_i0_i2 (.D(pc_5__N_35[2]), .SP(clk_c_enable_26), .CK(clk_c), 
            .Q(pc[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam pc_i0_i2.GSR = "ENABLED";
    FD1P3AX pc_i0_i1 (.D(pc_5__N_35[1]), .SP(clk_c_enable_26), .CK(clk_c), 
            .Q(pc[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam pc_i0_i1.GSR = "ENABLED";
    LUT4 div_28_i150_3_lut_rep_901_4_lut (.A(n46049), .B(n22715), .C(n46047), 
         .D(n23881), .Z(n46022)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (D))+!A (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_i150_3_lut_rep_901_4_lut.init = 16'h0df2;
    FD1S3IX states__i1 (.D(n3668[1]), .CK(clk_c), .CD(n22192), .Q(\states[1] )) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam states__i1.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut_adj_81 (.A(n396[7]), .B(n45917), .C(n45863), .D(n43750), 
         .Z(n23490)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(D)) */ ;
    defparam i1_2_lut_4_lut_adj_81.init = 16'h807f;
    LUT4 i15818_4_lut (.A(akku_o_c_4), .B(akku_o_8__N_67[4]), .C(n46276), 
         .D(data[4]), .Z(n22545)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(73[13] 82[22])
    defparam i15818_4_lut.init = 16'hc0c5;
    LUT4 n183_bdd_3_lut_4_lut (.A(n46049), .B(n22715), .C(n46037), .D(n46058), 
         .Z(n213)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (D))+!A (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam n183_bdd_3_lut_4_lut.init = 16'h0df2;
    LUT4 i1_4_lut_3_lut_rep_1150 (.A(akku_o_c_3), .B(akku_o_c_2), .C(akku_o_c_4), 
         .Z(n46271)) /* synthesis lut_function=(A (B (C))+!A !(B (C)+!B !(C))) */ ;
    defparam i1_4_lut_3_lut_rep_1150.init = 16'h9494;
    LUT4 i2_3_lut_4_lut_4_lut (.A(n3[2]), .B(n41242), .C(n3[1]), .D(n40849), 
         .Z(n40744)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_4_lut_4_lut.init = 16'h42bd;
    CCU2D div_28_add_187_9 (.A0(n22716), .B0(n46004), .C0(n231[7]), .D0(n212), 
          .A1(n22716), .B1(n46004), .C1(n231[8]), .D1(n211), .CIN(n40539), 
          .S0(n261[7]), .S1(n261[8]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_add_187_9.INIT0 = 16'h0e1f;
    defparam div_28_add_187_9.INIT1 = 16'h0e1f;
    defparam div_28_add_187_9.INJECT1_0 = "NO";
    defparam div_28_add_187_9.INJECT1_1 = "NO";
    LUT4 n338_bdd_3_lut_4_lut (.A(n45865), .B(n45872), .C(n541[4]), .D(n330[2]), 
         .Z(n45570)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C)+!B !(D)))) */ ;
    defparam n338_bdd_3_lut_4_lut.init = 16'h60f9;
    CCU2D div_28_add_187_7 (.A0(n22716), .B0(n46004), .C0(n231[5]), .D0(n46022), 
          .A1(n22716), .B1(n46004), .C1(n231[6]), .D1(n213), .CIN(n40538), 
          .COUT(n40539), .S0(n261[5]), .S1(n261[6]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_add_187_7.INIT0 = 16'h0e1f;
    defparam div_28_add_187_7.INIT1 = 16'h0e1f;
    defparam div_28_add_187_7.INJECT1_0 = "NO";
    defparam div_28_add_187_7.INJECT1_1 = "NO";
    CCU2D div_28_add_187_5 (.A0(n46029), .B0(n46155), .C0(n231[3]), .D0(n45991), 
          .A1(n22716), .B1(n46004), .C1(n231[4]), .D1(n215), .CIN(n40537), 
          .COUT(n40538), .S0(n261[3]), .S1(n261[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_add_187_5.INIT0 = 16'h0f66;
    defparam div_28_add_187_5.INIT1 = 16'h0e1f;
    defparam div_28_add_187_5.INJECT1_0 = "NO";
    defparam div_28_add_187_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_601_3_lut_4_lut_4_lut_4_lut (.A(n45730), .B(n45728), 
         .C(n45735), .D(n45724), .Z(n45722)) /* synthesis lut_function=(A (B+(C+(D)))+!A ((C+(D))+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_rep_601_3_lut_4_lut_4_lut_4_lut.init = 16'hfff9;
    LUT4 mux_181_i4_3_lut_4_lut (.A(n2203[5]), .B(n43670), .C(n46138), 
         .D(n45757), .Z(n825[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam mux_181_i4_3_lut_4_lut.init = 16'hf909;
    PFUMX i57 (.BLUT(n43557), .ALUT(n43532), .C0(akku_o_c_4), .Z(n31_adj_319));
    LUT4 i1_2_lut_rep_924_4_lut (.A(n46145), .B(n89_adj_320), .C(n46066), 
         .D(n46090), .Z(n46045)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_924_4_lut.init = 16'h2000;
    CCU2D add_277_3 (.A0(n999[0]), .B0(n999[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n999[1]), .B1(n999[5]), .C1(GND_net), .D1(GND_net), .CIN(n40422), 
          .COUT(n40423), .S0(n1012[1]), .S1(n1012[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_277_3.INIT0 = 16'h5999;
    defparam add_277_3.INIT1 = 16'h5999;
    defparam add_277_3.INJECT1_0 = "NO";
    defparam add_277_3.INJECT1_1 = "NO";
    CCU2D div_28_add_187_3 (.A0(akku_o_c_0), .B0(oprand[0]), .C0(n16[2]), 
          .D0(n16[1]), .A1(n46021), .B1(n22716), .C1(n231[2]), .D1(n217), 
          .CIN(n40536), .COUT(n40537), .S0(n261[1]), .S1(n261[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_add_187_3.INIT0 = 16'hfe10;
    defparam div_28_add_187_3.INIT1 = 16'hf1c0;
    defparam div_28_add_187_3.INJECT1_0 = "NO";
    defparam div_28_add_187_3.INJECT1_1 = "NO";
    LUT4 i5745_4_lut_3_lut (.A(n1324[5]), .B(n545[0]), .C(n1324[0]), .Z(n2)) /* synthesis lut_function=(A (B+(C))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5745_4_lut_3_lut.init = 16'he8e8;
    CCU2D div_28_add_187_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(akku_o_c_0), .B1(oprand[0]), .C1(n16[1]), 
          .D1(n16[0]), .COUT(n40536));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_add_187_1.INIT0 = 16'h0000;
    defparam div_28_add_187_1.INIT1 = 16'h01ef;
    defparam div_28_add_187_1.INJECT1_0 = "NO";
    defparam div_28_add_187_1.INJECT1_1 = "NO";
    LUT4 i2_3_lut_4_lut_4_lut_adj_82 (.A(n45794), .B(n45823), .C(n45790), 
         .D(n1687[5]), .Z(n40740)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D))+!B !(C (D)))) */ ;
    defparam i2_3_lut_4_lut_4_lut_adj_82.init = 16'hc933;
    LUT4 i31563_4_lut (.A(n23044), .B(n45822), .C(n21753), .D(n45892), 
         .Z(n38297)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i31563_4_lut.init = 16'h5455;
    LUT4 i2690_3_lut_4_lut_4_lut_4_lut (.A(n3[2]), .B(n41242), .C(n3[1]), 
         .D(n40849), .Z(n6_adj_321)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A !(B (C+!(D))+!B !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2690_3_lut_4_lut_4_lut_4_lut.init = 16'h40fd;
    LUT4 i2_2_lut_4_lut_3_lut (.A(akku_o_c_3), .B(akku_o_c_2), .C(akku_o_c_4), 
         .Z(n7_adj_322)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+(C))) */ ;
    defparam i2_2_lut_4_lut_3_lut.init = 16'hd6d6;
    CCU2D div_28_add_166_7 (.A0(n22715), .B0(n46049), .C0(n46028), .D0(n182), 
          .A1(n22715), .B1(n46049), .C1(n46020), .D1(n181), .CIN(n40534), 
          .S0(n231[7]), .S1(n231[8]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_add_166_7.INIT0 = 16'h0bf4;
    defparam div_28_add_166_7.INIT1 = 16'h0bf4;
    defparam div_28_add_166_7.INJECT1_0 = "NO";
    defparam div_28_add_166_7.INJECT1_1 = "NO";
    LUT4 div_39_i134_3_lut_rep_884_4_lut (.A(n46038), .B(n46050), .C(n169), 
         .D(n46039), .Z(n46005)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (C (D)+!C !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_i134_3_lut_rep_884_4_lut.init = 16'hf20d;
    LUT4 akku_o_c_3_bdd_4_lut_38331_4_lut (.A(akku_o_c_3), .B(akku_o_c_2), 
         .C(akku_o_c_4), .D(akku_o_c_1), .Z(n117_adj_323)) /* synthesis lut_function=(!((B (C (D)))+!A)) */ ;
    defparam akku_o_c_3_bdd_4_lut_38331_4_lut.init = 16'h2aaa;
    LUT4 i37283_4_lut (.A(n18[7]), .B(n44028), .C(n18[4]), .D(n43834), 
         .Z(n44177)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i37283_4_lut.init = 16'hfffe;
    LUT4 i37277_4_lut (.A(n221), .B(n44030), .C(n224), .D(n45970), .Z(n44171)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i37277_4_lut.init = 16'hfffe;
    CCU2D div_28_add_166_5 (.A0(n46022), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n46049), .B1(n46058), .C1(n201[6]), .D1(n22715), .CIN(n40533), 
          .COUT(n40534), .S0(n231[5]), .S1(n231[6]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_add_166_5.INIT0 = 16'h5555;
    defparam div_28_add_166_5.INIT1 = 16'h0f8d;
    defparam div_28_add_166_5.INJECT1_0 = "NO";
    defparam div_28_add_166_5.INJECT1_1 = "NO";
    CCU2D div_28_add_166_3 (.A0(n22715), .B0(n46057), .C0(n8_adj_310), 
          .D0(n46155), .A1(n46155), .B1(n46057), .C1(n22715), .D1(n41054), 
          .CIN(n40532), .COUT(n40533), .S0(n231[3]), .S1(n231[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_add_166_3.INIT0 = 16'hf4a0;
    defparam div_28_add_166_3.INIT1 = 16'h0cfe;
    defparam div_28_add_166_3.INJECT1_0 = "NO";
    defparam div_28_add_166_3.INJECT1_1 = "NO";
    LUT4 i37279_2_lut_rep_889_3_lut_4_lut (.A(n46061), .B(n46042), .C(n46062), 
         .Z(n46010)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i37279_2_lut_rep_889_3_lut_4_lut.init = 16'hf8f8;
    CCU2D div_28_add_166_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n46880), .B1(n46882), .C1(n16[3]), .D1(n16[2]), 
          .COUT(n40532), .S1(n231[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_add_166_1.INIT0 = 16'hF000;
    defparam div_28_add_166_1.INIT1 = 16'h01ef;
    defparam div_28_add_166_1.INJECT1_0 = "NO";
    defparam div_28_add_166_1.INJECT1_1 = "NO";
    CCU2D div_53_add_172_7 (.A0(n4_adj_325), .B0(n12), .C0(n45931), .D0(n191_adj_326), 
          .A1(n45946), .B1(n12), .C1(n45927), .D1(n45961), .CIN(n40530), 
          .S0(n20[7]), .S1(n20[8]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_add_172_7.INIT0 = 16'h0ff4;
    defparam div_53_add_172_7.INIT1 = 16'h0bf4;
    defparam div_53_add_172_7.INJECT1_0 = "NO";
    defparam div_53_add_172_7.INJECT1_1 = "NO";
    CCU2D div_53_add_172_5 (.A0(n12), .B0(n45953), .C0(n41038), .D0(n45946), 
          .A1(n45946), .B1(n12), .C1(n45945), .D1(n45954), .CIN(n40529), 
          .COUT(n40530), .S0(n20[5]), .S1(n20[6]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_add_172_5.INIT0 = 16'h0f8d;
    defparam div_53_add_172_5.INIT1 = 16'h0bf4;
    defparam div_53_add_172_5.INJECT1_0 = "NO";
    defparam div_53_add_172_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_879_3_lut_4_lut_4_lut (.A(n46061), .B(n46042), .C(n46062), 
         .Z(n46000)) /* synthesis lut_function=(A (B+!(C))+!A (B (C)+!B !(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_rep_879_3_lut_4_lut_4_lut.init = 16'hcbcb;
    CCU2D div_53_add_172_3 (.A0(n45946), .B0(n43883), .C0(n8_adj_331), 
          .D0(n45975), .A1(n12), .B1(n45952), .C1(n45943), .D1(n45946), 
          .CIN(n40528), .COUT(n40529), .S0(n20[3]), .S1(n20[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_add_172_3.INIT0 = 16'hf4a0;
    defparam div_53_add_172_3.INIT1 = 16'hf072;
    defparam div_53_add_172_3.INJECT1_0 = "NO";
    defparam div_53_add_172_3.INJECT1_1 = "NO";
    CCU2D div_53_add_172_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n22712), .B1(n45965), .C1(n46123), .D1(n45944), 
          .COUT(n40528), .S1(n20[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_add_172_1.INIT0 = 16'hF000;
    defparam div_53_add_172_1.INIT1 = 16'h04f4;
    defparam div_53_add_172_1.INJECT1_0 = "NO";
    defparam div_53_add_172_1.INJECT1_1 = "NO";
    CCU2D div_53_add_193_9 (.A0(n22673), .B0(n45922), .C0(n20[7]), .D0(n221_adj_333), 
          .A1(n22673), .B1(n45922), .C1(n20[8]), .D1(n220), .CIN(n40526), 
          .S0(n270[7]), .S1(n270[8]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_add_193_9.INIT0 = 16'h0e1f;
    defparam div_53_add_193_9.INIT1 = 16'h0e1f;
    defparam div_53_add_193_9.INJECT1_0 = "NO";
    defparam div_53_add_193_9.INJECT1_1 = "NO";
    PFUMX i38439 (.BLUT(n46296), .ALUT(n46297), .C0(n46873), .Z(n59));
    CCU2D div_53_add_193_7 (.A0(n22673), .B0(n45922), .C0(n20[5]), .D0(n223), 
          .A1(n22673), .B1(n45922), .C1(n20[6]), .D1(n222_adj_334), 
          .CIN(n40525), .COUT(n40526), .S0(n270[5]), .S1(n270[6]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_add_193_7.INIT0 = 16'h0e1f;
    defparam div_53_add_193_7.INIT1 = 16'h0e1f;
    defparam div_53_add_193_7.INJECT1_0 = "NO";
    defparam div_53_add_193_7.INJECT1_1 = "NO";
    LUT4 div_46_i133_3_lut_4_lut_3_lut_4_lut (.A(n46061), .B(n46042), .C(n46062), 
         .Z(n191_adj_335)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_46_i133_3_lut_4_lut_3_lut_4_lut.init = 16'h8080;
    CCU2D div_53_add_193_5 (.A0(n45932), .B0(n45975), .C0(n20[3]), .D0(n45916), 
          .A1(n22673), .B1(n45922), .C1(n20[4]), .D1(n45925), .CIN(n40524), 
          .COUT(n40525), .S0(n270[3]), .S1(n270[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_add_193_5.INIT0 = 16'hf099;
    defparam div_53_add_193_5.INIT1 = 16'h0e1f;
    defparam div_53_add_193_5.INJECT1_0 = "NO";
    defparam div_53_add_193_5.INJECT1_1 = "NO";
    LUT4 i33208_2_lut_rep_1102_3_lut (.A(akku_o_c_2), .B(akku_o_c_1), .C(akku_o_c_3), 
         .Z(n46223)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i33208_2_lut_rep_1102_3_lut.init = 16'hf8f8;
    CCU2D div_53_add_193_3 (.A0(n43353), .B0(n45937), .C0(n46123), .D0(n107), 
          .A1(n22035), .B1(n22673), .C1(n20[2]), .D1(n73_adj_336), .CIN(n40523), 
          .COUT(n40524), .S0(n270[1]), .S1(n270[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_add_193_3.INIT0 = 16'hfe0e;
    defparam div_53_add_193_3.INIT1 = 16'hf1c0;
    defparam div_53_add_193_3.INJECT1_0 = "NO";
    defparam div_53_add_193_3.INJECT1_1 = "NO";
    CCU2D div_53_add_193_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n43333), .B1(n30878), .C1(n46123), .D1(n108), 
          .COUT(n40523));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_add_193_1.INIT0 = 16'h0000;
    defparam div_53_add_193_1.INIT1 = 16'h01f1;
    defparam div_53_add_193_1.INJECT1_0 = "NO";
    defparam div_53_add_193_1.INJECT1_1 = "NO";
    LUT4 div_46_i134_3_lut_rep_876_4_lut_4_lut (.A(n46061), .B(n46042), 
         .C(n46062), .Z(n45997)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_46_i134_3_lut_rep_876_4_lut_4_lut.init = 16'h6262;
    CCU2D add_277_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n30783), .B1(n16[8]), .C1(n46196), .D1(n462[4]), .COUT(n40422), 
          .S1(n1012[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_277_1.INIT0 = 16'hF000;
    defparam add_277_1.INIT1 = 16'h07f7;
    defparam add_277_1.INJECT1_0 = "NO";
    defparam add_277_1.INJECT1_1 = "NO";
    LUT4 i33696_2_lut_rep_1052_3_lut_4_lut_4_lut (.A(akku_o_c_2), .B(akku_o_c_1), 
         .C(akku_o_c_4), .D(akku_o_c_3), .Z(n46173)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B (C (D))+!B !(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i33696_2_lut_rep_1052_3_lut_4_lut_4_lut.init = 16'h3c4c;
    CCU2D add_1769_9 (.A0(akku_o_c_7), .B0(data_7__N_89[7]), .C0(data_7__N_102), 
          .D0(n46197), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n40522), .S0(akku_o_8__N_67[7]), .S1(akku_o_8__N_67[8]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(74[39:69])
    defparam add_1769_9.INIT0 = 16'h556a;
    defparam add_1769_9.INIT1 = 16'h0000;
    defparam add_1769_9.INJECT1_0 = "NO";
    defparam add_1769_9.INJECT1_1 = "NO";
    CCU2D add_1769_7 (.A0(akku_o_c_5), .B0(data_7__N_89[5]), .C0(data_7__N_102), 
          .D0(n46199), .A1(akku_o_c_6), .B1(data_7__N_89[6]), .C1(data_7__N_102), 
          .D1(n46198), .CIN(n40521), .COUT(n40522), .S0(akku_o_8__N_67[5]), 
          .S1(akku_o_8__N_67[6]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(74[39:69])
    defparam add_1769_7.INIT0 = 16'h556a;
    defparam add_1769_7.INIT1 = 16'h556a;
    defparam add_1769_7.INJECT1_0 = "NO";
    defparam add_1769_7.INJECT1_1 = "NO";
    CCU2D add_1769_5 (.A0(akku_o_c_3), .B0(data_7__N_89[3]), .C0(data_7__N_102), 
          .D0(n46200), .A1(akku_o_c_4), .B1(data_7__N_89[4]), .C1(data_7__N_102), 
          .D1(n46175), .CIN(n40520), .COUT(n40521), .S0(akku_o_8__N_67[3]), 
          .S1(akku_o_8__N_67[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(74[39:69])
    defparam add_1769_5.INIT0 = 16'h556a;
    defparam add_1769_5.INIT1 = 16'h556a;
    defparam add_1769_5.INJECT1_0 = "NO";
    defparam add_1769_5.INJECT1_1 = "NO";
    CCU2D add_1769_3 (.A0(akku_o_c_1), .B0(data_7__N_89[1]), .C0(data_7__N_102), 
          .D0(n46202), .A1(akku_o_c_2), .B1(data_7__N_89[2]), .C1(data_7__N_102), 
          .D1(n46201), .CIN(n40519), .COUT(n40520), .S0(akku_o_8__N_67[1]), 
          .S1(akku_o_8__N_67[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(74[39:69])
    defparam add_1769_3.INIT0 = 16'h556a;
    defparam add_1769_3.INIT1 = 16'h556a;
    defparam add_1769_3.INJECT1_0 = "NO";
    defparam add_1769_3.INJECT1_1 = "NO";
    LUT4 i37285_4_lut (.A(n30723), .B(n44099), .C(n44026), .D(n270_adj_514[2]), 
         .Z(n44179)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i37285_4_lut.init = 16'hfefc;
    CCU2D add_1769_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(akku_o_c_0), .B1(data_7__N_89[0]), .C1(data_7__N_102), .D1(n46181), 
          .COUT(n40519), .S1(n4247[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(74[39:69])
    defparam add_1769_1.INIT0 = 16'hF000;
    defparam add_1769_1.INIT1 = 16'h556a;
    defparam add_1769_1.INJECT1_0 = "NO";
    defparam add_1769_1.INJECT1_1 = "NO";
    CCU2D add_613_7 (.A0(n2616[4]), .B0(n2616[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40518), 
          .S0(n2629[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_613_7.INIT0 = 16'h5999;
    defparam add_613_7.INIT1 = 16'h0000;
    defparam add_613_7.INJECT1_0 = "NO";
    defparam add_613_7.INJECT1_1 = "NO";
    CCU2D add_613_5 (.A0(n2616[2]), .B0(n2616[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2616[3]), .B1(n2616[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40517), .COUT(n40518), .S0(n2629[3]), .S1(n2629[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_613_5.INIT0 = 16'h5666;
    defparam add_613_5.INIT1 = 16'h5666;
    defparam add_613_5.INJECT1_0 = "NO";
    defparam add_613_5.INJECT1_1 = "NO";
    CCU2D add_613_3 (.A0(n2616[0]), .B0(n2616[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2616[1]), .B1(n2616[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40516), .COUT(n40517), .S0(n2629[1]), .S1(n2629[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_613_3.INIT0 = 16'h5999;
    defparam add_613_3.INIT1 = 16'h5666;
    defparam add_613_3.INJECT1_0 = "NO";
    defparam add_613_3.INJECT1_1 = "NO";
    LUT4 mux_33_i7_4_lut (.A(n16[8]), .B(n112[6]), .C(n46207), .D(n46120), 
         .Z(n102)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_33_i7_4_lut.init = 16'hcac0;
    LUT4 i1_2_lut_rep_919_4_lut (.A(n46136), .B(n46060), .C(n22585), .D(n46104), 
         .Z(n46040)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_919_4_lut.init = 16'h8000;
    LUT4 i31995_2_lut_rep_916_3_lut_4_lut (.A(n46143), .B(n46852), .C(n23881), 
         .D(n46155), .Z(n46037)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(B (C)+!B !((D)+!C))) */ ;
    defparam i31995_2_lut_rep_916_3_lut_4_lut.init = 16'h9f0f;
    LUT4 i37292_3_lut (.A(n45942), .B(n44181), .C(n30723), .Z(n44187)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i37292_3_lut.init = 16'hecec;
    LUT4 i1_3_lut_4_lut (.A(n396[7]), .B(n45917), .C(n45863), .D(n45849), 
         .Z(n22969)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf08f;
    LUT4 i1_2_lut_rep_923_4_lut (.A(n46136), .B(n46060), .C(n22585), .D(n46111), 
         .Z(n46044)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_923_4_lut.init = 16'h8000;
    LUT4 i15802_4_lut (.A(akku_o_8__N_50[1]), .B(n43707), .C(n46854), 
         .D(n3622), .Z(n22529)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(73[13] 82[22])
    defparam i15802_4_lut.init = 16'hca0a;
    PFUMX i38192 (.BLUT(n45285), .ALUT(n45284), .C0(n86), .Z(n45286));
    CCU2D add_613_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n8_adj_338), .B1(n46209), .C1(n43349), .D1(n860[1]), .COUT(n40516), 
          .S1(n2629[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_613_1.INIT0 = 16'hF000;
    defparam add_613_1.INIT1 = 16'h01ff;
    defparam add_613_1.INJECT1_0 = "NO";
    defparam add_613_1.INJECT1_1 = "NO";
    CCU2D add_611_7 (.A0(n2603[4]), .B0(n2603[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40515), 
          .S0(n2616[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_611_7.INIT0 = 16'h5999;
    defparam add_611_7.INIT1 = 16'h0000;
    defparam add_611_7.INJECT1_0 = "NO";
    defparam add_611_7.INJECT1_1 = "NO";
    CCU2D add_611_5 (.A0(n2603[2]), .B0(n2603[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2603[3]), .B1(n2603[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40514), .COUT(n40515), .S0(n2616[3]), .S1(n2616[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_611_5.INIT0 = 16'h5666;
    defparam add_611_5.INIT1 = 16'h5666;
    defparam add_611_5.INJECT1_0 = "NO";
    defparam add_611_5.INJECT1_1 = "NO";
    CCU2D add_611_3 (.A0(n2603[0]), .B0(n2603[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2603[1]), .B1(n2603[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40513), .COUT(n40514), .S0(n2616[1]), .S1(n2616[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_611_3.INIT0 = 16'h5999;
    defparam add_611_3.INIT1 = 16'h5666;
    defparam add_611_3.INJECT1_0 = "NO";
    defparam add_611_3.INJECT1_1 = "NO";
    CCU2D add_611_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n43712), .B1(n45731), .C1(n46157), .D1(n45738), .COUT(n40513), 
          .S1(n2616[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_611_1.INIT0 = 16'hF000;
    defparam add_611_1.INIT1 = 16'h09f9;
    defparam add_611_1.INJECT1_0 = "NO";
    defparam add_611_1.INJECT1_1 = "NO";
    CCU2D add_609_7 (.A0(n2590[4]), .B0(n2590[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40512), 
          .S0(n2603[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_609_7.INIT0 = 16'h5999;
    defparam add_609_7.INIT1 = 16'h0000;
    defparam add_609_7.INJECT1_0 = "NO";
    defparam add_609_7.INJECT1_1 = "NO";
    CCU2D add_609_5 (.A0(n2590[2]), .B0(n2590[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2590[3]), .B1(n2590[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40511), .COUT(n40512), .S0(n2603[3]), .S1(n2603[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_609_5.INIT0 = 16'h5666;
    defparam add_609_5.INIT1 = 16'h5666;
    defparam add_609_5.INJECT1_0 = "NO";
    defparam add_609_5.INJECT1_1 = "NO";
    CCU2D add_609_3 (.A0(n2590[0]), .B0(n2590[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2590[1]), .B1(n2590[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40510), .COUT(n40511), .S0(n2603[1]), .S1(n2603[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_609_3.INIT0 = 16'h5999;
    defparam add_609_3.INIT1 = 16'h5666;
    defparam add_609_3.INJECT1_0 = "NO";
    defparam add_609_3.INJECT1_1 = "NO";
    CCU2D add_609_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n43673), .B1(n7_adj_339), .C1(n46157), .D1(n45743), .COUT(n40510), 
          .S1(n2603[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_609_1.INIT0 = 16'hF000;
    defparam add_609_1.INIT1 = 16'h06f6;
    defparam add_609_1.INJECT1_0 = "NO";
    defparam add_609_1.INJECT1_1 = "NO";
    CCU2D add_607_7 (.A0(n2577[4]), .B0(n2577[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40509), 
          .S0(n2590[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_607_7.INIT0 = 16'h5999;
    defparam add_607_7.INIT1 = 16'h0000;
    defparam add_607_7.INJECT1_0 = "NO";
    defparam add_607_7.INJECT1_1 = "NO";
    CCU2D add_607_5 (.A0(n2577[2]), .B0(n2577[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2577[3]), .B1(n2577[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40508), .COUT(n40509), .S0(n2590[3]), .S1(n2590[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_607_5.INIT0 = 16'h5666;
    defparam add_607_5.INIT1 = 16'h5666;
    defparam add_607_5.INJECT1_0 = "NO";
    defparam add_607_5.INJECT1_1 = "NO";
    LUT4 mux_47_i7_4_lut_rep_1165 (.A(n46096), .B(n46083), .C(n46123), 
         .D(n46097), .Z(n46851)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_47_i7_4_lut_rep_1165.init = 16'hcac0;
    LUT4 i1_2_lut_rep_741_4_lut (.A(n45866), .B(n3[3]), .C(n37_adj_340), 
         .D(n45872), .Z(n45862)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(B (D)+!B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_741_4_lut.init = 16'ha35c;
    LUT4 mux_72_i5_3_lut (.A(n45908), .B(n45915), .C(n43592), .Z(n3[4])) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_72_i5_3_lut.init = 16'h5c5c;
    LUT4 rem_87_i85_3_lut_4_lut_4_lut_4_lut_3_lut_4_lut (.A(oprand[1]), .B(n46876), 
         .C(n46873), .D(oprand[3]), .Z(n118_adj_306)) /* synthesis lut_function=(A (B)+!A !((C (D))+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(20[15:21])
    defparam rem_87_i85_3_lut_4_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h8ccc;
    LUT4 i4995_3_lut_4_lut_4_lut (.A(n2203[5]), .B(n45751), .C(n6_adj_341), 
         .D(n43670), .Z(n8_adj_342)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B ((D)+!C)+!B !(C+!(D)))) */ ;
    defparam i4995_3_lut_4_lut_4_lut.init = 16'hb8d1;
    LUT4 mux_79_i2_3_lut_rep_724_4_lut (.A(n449[4]), .B(n3[1]), .C(n39), 
         .D(n51), .Z(n45845)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_79_i2_3_lut_rep_724_4_lut.init = 16'h5ccc;
    LUT4 mux_40_i5_3_lut_rep_888_4_lut (.A(n169), .B(n46050), .C(n31), 
         .D(n43_adj_299), .Z(n46009)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_40_i5_3_lut_rep_888_4_lut.init = 16'h5ccc;
    LUT4 mux_93_i4_3_lut_rep_715_4_lut (.A(n41291), .B(n45848), .C(n39_adj_343), 
         .D(n51_adj_344), .Z(n45836)) /* synthesis lut_function=(A (B+(C (D)))+!A !((C (D))+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_93_i4_3_lut_rep_715_4_lut.init = 16'haccc;
    LUT4 mux_40_i1_3_lut_4_lut (.A(n55), .B(n168), .C(n31), .D(n43_adj_299), 
         .Z(n108)) /* synthesis lut_function=(A (B+(C (D)))+!A !((C (D))+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_40_i1_3_lut_4_lut.init = 16'haccc;
    LUT4 mux_93_i3_3_lut_rep_695_4_lut (.A(n45819), .B(n363[2]), .C(n39_adj_343), 
         .D(n51_adj_344), .Z(n45816)) /* synthesis lut_function=(A (B+(C (D)))+!A !((C (D))+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_93_i3_3_lut_rep_695_4_lut.init = 16'haccc;
    LUT4 mux_188_i4_3_lut_rep_622_4_lut (.A(n2345[5]), .B(n825[3]), .C(n45390), 
         .D(n59), .Z(n45743)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_188_i4_3_lut_rep_622_4_lut.init = 16'h5ccc;
    LUT4 mux_107_i6_3_lut_4_lut (.A(n866[4]), .B(n45859), .C(n39_adj_313), 
         .D(n51_adj_345), .Z(n462[5])) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_107_i6_3_lut_4_lut.init = 16'h5ccc;
    LUT4 i1_2_lut_rep_745 (.A(n43720), .B(n43729), .Z(n45866)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_rep_745.init = 16'h6666;
    LUT4 mux_188_i3_3_lut_rep_617_4_lut (.A(n2358[5]), .B(n825[2]), .C(n45390), 
         .D(n59), .Z(n45738)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_188_i3_3_lut_rep_617_4_lut.init = 16'h5ccc;
    LUT4 i14917_3_lut_rep_743_4_lut (.A(n43720), .B(n43729), .C(n3[2]), 
         .D(n3[3]), .Z(n45864)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (B (D)+!B ((D)+!C)))) */ ;
    defparam i14917_3_lut_rep_743_4_lut.init = 16'h00f6;
    LUT4 mux_188_i2_3_lut_4_lut (.A(n2371[5]), .B(n825[1]), .C(n45390), 
         .D(n59), .Z(n860[1])) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_188_i2_3_lut_4_lut.init = 16'h5ccc;
    LUT4 i1_2_lut_rep_1008_3_lut_4_lut (.A(n46177), .B(n43349), .C(n45390), 
         .D(n59), .Z(n46129)) /* synthesis lut_function=(!(A (C (D))+!A ((C (D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_2_lut_rep_1008_3_lut_4_lut.init = 16'h0eee;
    CCU2D add_607_3 (.A0(n2577[0]), .B0(n2577[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2577[1]), .B1(n2577[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40507), .COUT(n40508), .S0(n2590[1]), .S1(n2590[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_607_3.INIT0 = 16'h5999;
    defparam add_607_3.INIT1 = 16'h5666;
    defparam add_607_3.INJECT1_0 = "NO";
    defparam add_607_3.INJECT1_1 = "NO";
    LUT4 i4852_2_lut_rep_895_4_lut (.A(n46090), .B(n46041), .C(n43581), 
         .D(n825[7]), .Z(n46016)) /* synthesis lut_function=(!(A (B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i4852_2_lut_rep_895_4_lut.init = 16'h7fff;
    LUT4 mux_107_i2_3_lut_4_lut (.A(n910[4]), .B(n429[1]), .C(n39_adj_313), 
         .D(n51_adj_345), .Z(n462[1])) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_107_i2_3_lut_4_lut.init = 16'h5ccc;
    LUT4 mux_40_i2_3_lut_4_lut (.A(n146[1]), .B(n257), .C(n31), .D(n43_adj_299), 
         .Z(n107)) /* synthesis lut_function=(A (B+(C (D)))+!A !((C (D))+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_40_i2_3_lut_4_lut.init = 16'haccc;
    LUT4 mux_54_i2_3_lut_4_lut (.A(n208[1]), .B(n107_adj_346), .C(n45287), 
         .D(n45286), .Z(n218[1])) /* synthesis lut_function=(A (B+(C (D)))+!A !((C (D))+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_54_i2_3_lut_4_lut.init = 16'haccc;
    LUT4 n44042_bdd_4_lut (.A(n46171), .B(n46240), .C(n46261), .D(n46873), 
         .Z(n45481)) /* synthesis lut_function=(A+!(B (C+!(D)))) */ ;
    defparam n44042_bdd_4_lut.init = 16'hbfbb;
    LUT4 mux_107_i3_3_lut_4_lut (.A(n45807), .B(n429[2]), .C(n39_adj_313), 
         .D(n51_adj_345), .Z(n462[2])) /* synthesis lut_function=(A (B+(C (D)))+!A !((C (D))+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_107_i3_3_lut_4_lut.init = 16'haccc;
    LUT4 mux_79_i6_3_lut_rep_803_4_lut (.A(n45929), .B(n45940), .C(n39), 
         .D(n51), .Z(n45924)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_79_i6_3_lut_rep_803_4_lut.init = 16'h5ccc;
    LUT4 i23732_4_lut (.A(n40781), .B(n19), .C(n685[0]), .D(n89), .Z(n755[0])) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i23732_4_lut.init = 16'h88c0;
    LUT4 i23862_2_lut_rep_793_3_lut_4_lut (.A(n45923), .B(n39_adj_343), 
         .C(n51_adj_344), .D(n15_adj_316), .Z(n45914)) /* synthesis lut_function=(!((B (C+!(D))+!B !(D))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i23862_2_lut_rep_793_3_lut_4_lut.init = 16'h2a00;
    LUT4 akku_o_c_1_bdd_4_lut_4_lut (.A(akku_o_c_1), .B(akku_o_c_2), .C(akku_o_c_4), 
         .D(akku_o_c_3), .Z(n44162)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A (B+(D))) */ ;
    defparam akku_o_c_1_bdd_4_lut_4_lut.init = 16'hff6e;
    LUT4 mux_167_i7_4_lut (.A(n45788), .B(n89), .C(n19), .D(n45892), 
         .Z(n755[6])) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_167_i7_4_lut.init = 16'h3a0a;
    LUT4 i37009_2_lut_rep_993_3_lut (.A(n43592), .B(n39), .C(n51), .Z(n46114)) /* synthesis lut_function=(A+(B (C))) */ ;
    defparam i37009_2_lut_rep_993_3_lut.init = 16'heaea;
    LUT4 mux_79_i3_3_lut_4_lut (.A(n41242), .B(n3[2]), .C(n39), .D(n51), 
         .Z(n330[2])) /* synthesis lut_function=(A (B+(C (D)))+!A !((C (D))+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_79_i3_3_lut_4_lut.init = 16'haccc;
    LUT4 i1_2_lut_3_lut_4_lut_adj_83 (.A(n45762), .B(n45754), .C(n43709), 
         .D(n2203[5]), .Z(n43710)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_83.init = 16'h6996;
    LUT4 mux_100_i4_3_lut_4_lut (.A(n43695), .B(n43750), .C(n45836), .D(n15_adj_316), 
         .Z(n429[3])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_100_i4_3_lut_4_lut.init = 16'hf099;
    LUT4 i2_3_lut_4_lut_adj_84 (.A(n43720), .B(n43729), .C(n22894), .D(n41385), 
         .Z(n449[4])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i2_3_lut_4_lut_adj_84.init = 16'h9669;
    CCU2D add_275_7 (.A0(VCC_net), .B0(n45900), .C0(n475[8]), .D0(n46035), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40421), 
          .S0(n999[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_275_7.INIT0 = 16'haaa9;
    defparam add_275_7.INIT1 = 16'h0000;
    defparam add_275_7.INJECT1_0 = "NO";
    defparam add_275_7.INJECT1_1 = "NO";
    LUT4 i2_4_lut (.A(n46409), .B(n3[8]), .C(n45933), .D(n6383), .Z(n43720)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i2_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_977_3_lut_4_lut (.A(n39_adj_343), .B(n51_adj_344), 
         .C(n46110), .D(n15_adj_316), .Z(n46098)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_977_3_lut_4_lut.init = 16'h7000;
    LUT4 mux_188_i5_3_lut_rep_637_4_lut (.A(n2332[5]), .B(n825[4]), .C(n45390), 
         .D(n59), .Z(n45758)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_188_i5_3_lut_rep_637_4_lut.init = 16'h5ccc;
    LUT4 i2_3_lut_4_lut_adj_85 (.A(n43720), .B(n43729), .C(n3[3]), .D(n3[2]), 
         .Z(n40849)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i2_3_lut_4_lut_adj_85.init = 16'h6996;
    LUT4 i2_4_lut_then_4_lut (.A(n2098[5]), .B(n2098[4]), .C(n2098[2]), 
         .D(n4_adj_347), .Z(n46281)) /* synthesis lut_function=(A (B)+!A !(B (C (D))+!B !(C (D)))) */ ;
    defparam i2_4_lut_then_4_lut.init = 16'h9ccc;
    LUT4 i5828_2_lut_4_lut (.A(n910[4]), .B(n429[1]), .C(n429[0]), .D(n4_adj_348), 
         .Z(n21933)) /* synthesis lut_function=(A+!(B+((D)+!C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5828_2_lut_4_lut.init = 16'haaba;
    LUT4 mux_79_i4_3_lut_rep_744_4_lut (.A(n43720), .B(n43729), .C(n37_adj_340), 
         .D(n3[3]), .Z(n45865)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;
    defparam mux_79_i4_3_lut_rep_744_4_lut.init = 16'h9f90;
    LUT4 i5827_2_lut_4_lut (.A(n910[4]), .B(n429[1]), .C(n429[0]), .D(n4_adj_348), 
         .Z(n9938)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5827_2_lut_4_lut.init = 16'haaa2;
    LUT4 i38071_4_lut_4_lut (.A(n44713), .B(n45732), .C(n45726), .D(n2734[3]), 
         .Z(n44699)) /* synthesis lut_function=(A (B (C (D))+!B !(D))+!A (B (D)+!B !(C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i38071_4_lut_4_lut.init = 16'hc533;
    LUT4 i3_4_lut_4_lut_adj_86 (.A(n46179), .B(n46875), .C(n46873), .D(n14), 
         .Z(n19)) /* synthesis lut_function=(A+(B ((D)+!C)+!B (C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    defparam i3_4_lut_4_lut_adj_86.init = 16'hffbe;
    LUT4 i5689_4_lut (.A(n1855[2]), .B(n2_adj_349), .C(n1855[5]), .D(n1855[1]), 
         .Z(n6_adj_350)) /* synthesis lut_function=(A (B+((D)+!C))+!A !((C+!(D))+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5689_4_lut.init = 16'hae8a;
    LUT4 i1_2_lut_3_lut_adj_87 (.A(n45762), .B(n45754), .C(n6_adj_341), 
         .Z(n4_adj_351)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i1_2_lut_3_lut_adj_87.init = 16'h9696;
    LUT4 i1_2_lut_rep_746 (.A(n46848), .B(n43759), .Z(n45867)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_rep_746.init = 16'h6666;
    LUT4 n935_bdd_4_lut (.A(n46845), .B(n45771), .C(n45749), .Z(n2734[3])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;
    defparam n935_bdd_4_lut.init = 16'h6c6c;
    CCU2D add_607_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n43349), .B1(n2476[5]), .C1(n46177), .D1(n45758), .COUT(n40507), 
          .S1(n2590[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_607_1.INIT0 = 16'hF000;
    defparam add_607_1.INIT1 = 16'h04fe;
    defparam add_607_1.INJECT1_0 = "NO";
    defparam add_607_1.INJECT1_1 = "NO";
    LUT4 i24460_4_lut_then_4_lut (.A(oprand[2]), .B(oprand[3]), .C(oprand[1]), 
         .D(oprand[4]), .Z(n46316)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;
    defparam i24460_4_lut_then_4_lut.init = 16'h7f80;
    LUT4 i24460_4_lut_else_4_lut (.A(oprand[2]), .B(oprand[3]), .C(oprand[1]), 
         .D(oprand[4]), .Z(n46315)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(D))) */ ;
    defparam i24460_4_lut_else_4_lut.init = 16'h7f00;
    LUT4 n117_bdd_4_lut_4_lut (.A(oprand[1]), .B(n46876), .C(n46875), 
         .D(n46873), .Z(n43941)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B+(C))) */ ;
    defparam n117_bdd_4_lut_4_lut.init = 16'hf6fe;
    LUT4 i7486_2_lut_rep_857_4_lut_else_4_lut_4_lut_4_lut (.A(n46096), .B(n46083), 
         .C(n46123), .D(n46097), .Z(n46850)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i7486_2_lut_rep_857_4_lut_else_4_lut_4_lut_4_lut.init = 16'h7000;
    LUT4 n1701_bdd_4_lut (.A(n45782), .B(n650[1]), .C(n45784), .D(n650[2]), 
         .Z(n45489)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A !(B ((D)+!C)+!B !(C)))) */ ;
    defparam n1701_bdd_4_lut.init = 16'h4fad;
    LUT4 mux_72_i3_3_lut_4_lut (.A(n46848), .B(n43759), .C(n43592), .D(n21[2]), 
         .Z(n3[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;
    defparam mux_72_i3_3_lut_4_lut.init = 16'h9f90;
    LUT4 i23731_4_lut (.A(n46406), .B(n46137), .C(n615[0]), .D(n89_adj_303), 
         .Z(n685[0])) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i23731_4_lut.init = 16'h88c0;
    LUT4 i2_2_lut_rep_935_4_lut (.A(n46851), .B(n46071), .C(n29_adj_353), 
         .D(n46179), .Z(n46056)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))) */ ;
    defparam i2_2_lut_rep_935_4_lut.init = 16'h8a00;
    LUT4 i1_4_lut_adj_88 (.A(n45694), .B(n46249), .C(akku_o_c_2), .D(n83), 
         .Z(n43564)) /* synthesis lut_function=(!(A (B)+!A (B+(C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_4_lut_adj_88.init = 16'h2322;
    LUT4 oprand_1__bdd_4_lut_38523 (.A(oprand[1]), .B(oprand[4]), .C(oprand[3]), 
         .D(n46876), .Z(n46318)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam oprand_1__bdd_4_lut_38523.init = 16'h18f0;
    LUT4 rem_61_i84_3_lut_4_lut_4_lut (.A(akku_o_c_3), .B(akku_o_c_2), .C(akku_o_c_1), 
         .D(akku_o_c_4), .Z(n117_adj_354)) /* synthesis lut_function=(A (B+(C+!(D)))) */ ;
    defparam rem_61_i84_3_lut_4_lut_4_lut.init = 16'ha8aa;
    LUT4 i24456_4_lut_then_4_lut (.A(akku_o_c_3), .B(akku_o_c_2), .C(akku_o_c_4), 
         .D(akku_o_c_1), .Z(n46320)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i24456_4_lut_then_4_lut.init = 16'h78f0;
    LUT4 i24456_4_lut_else_4_lut (.A(akku_o_c_3), .B(akku_o_c_2), .C(akku_o_c_4), 
         .D(akku_o_c_1), .Z(n46319)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;
    defparam i24456_4_lut_else_4_lut.init = 16'h70f0;
    LUT4 i133_then_4_lut (.A(oprand[2]), .B(oprand[0]), .C(oprand[4]), 
         .D(oprand[3]), .Z(n46323)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i133_then_4_lut.init = 16'h0040;
    LUT4 i133_else_4_lut (.A(oprand[2]), .B(oprand[0]), .C(oprand[3]), 
         .Z(n46322)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i133_else_4_lut.init = 16'h0101;
    CCU2D add_605_7 (.A0(n43991), .B0(n6_adj_355), .C0(n2662), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40506), 
          .S0(n2577[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_605_7.INIT0 = 16'he1e1;
    defparam add_605_7.INIT1 = 16'h0000;
    defparam add_605_7.INJECT1_0 = "NO";
    defparam add_605_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_89 (.A(n46090), .B(n46041), .C(n43581), .D(n46129), 
         .Z(n895[8])) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_4_lut_adj_89.init = 16'h8000;
    LUT4 i1_2_lut_4_lut_adj_90 (.A(n46128), .B(n45_adj_356), .C(n46074), 
         .D(n46090), .Z(n545[8])) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_4_lut_adj_90.init = 16'h2000;
    LUT4 i5911_2_lut_4_lut_4_lut (.A(n45902), .B(n40960), .C(n231_adj_515[0]), 
         .D(n4_adj_357), .Z(n10022)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5911_2_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 mux_65_i6_3_lut (.A(n22855), .B(n45987), .C(n37_adj_318), .Z(n293[1])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_65_i6_3_lut.init = 16'hacac;
    LUT4 i5912_2_lut_4_lut_4_lut (.A(n45902), .B(n40960), .C(n231_adj_515[0]), 
         .D(n4_adj_357), .Z(n21951)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5912_2_lut_4_lut_4_lut.init = 16'hfffd;
    LUT4 i15789_2_lut_rep_947_3_lut_4_lut_4_lut (.A(n46096), .B(n46083), 
         .C(n46123), .D(n46097), .Z(n46068)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A !(B (C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i15789_2_lut_rep_947_3_lut_4_lut_4_lut.init = 16'h4ac0;
    LUT4 i1_4_lut_adj_91 (.A(n46215), .B(n109), .C(n43606), .D(n40006), 
         .Z(n89)) /* synthesis lut_function=(A (B ((D)+!C))+!A !((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_4_lut_adj_91.init = 16'h8c0c;
    LUT4 i1_4_lut_adj_92 (.A(n46403), .B(n46385), .C(n46379), .D(n46873), 
         .Z(n109)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_4_lut_adj_92.init = 16'h40c0;
    LUT4 i132_then_4_lut (.A(akku_o_c_3), .B(akku_o_c_0), .C(akku_o_c_4), 
         .D(akku_o_c_2), .Z(n46329)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i132_then_4_lut.init = 16'h0040;
    LUT4 i2_3_lut_4_lut_4_lut_adj_93 (.A(n45869), .B(n45923), .C(n45856), 
         .D(n43686), .Z(n640[2])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;
    defparam i2_3_lut_4_lut_4_lut_adj_93.init = 16'h6c36;
    LUT4 i1_4_lut_rep_1166 (.A(n46088), .B(n12_adj_358), .C(n152), .Z(n46852)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i1_4_lut_rep_1166.init = 16'h0404;
    LUT4 i1_4_lut_then_4_lut (.A(oprand[3]), .B(oprand[2]), .C(oprand[1]), 
         .D(n6_adj_359), .Z(n46332)) /* synthesis lut_function=(A (B (C (D)))+!A !(B (C))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h9515;
    LUT4 i1_4_lut_else_4_lut (.A(oprand[3]), .B(n6_adj_359), .Z(n46331)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_927_3_lut_4_lut (.A(n15_adj_316), .B(n46075), .C(n46136), 
         .D(n37), .Z(n46048)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_927_3_lut_4_lut.init = 16'h0080;
    LUT4 i3049_3_lut_rep_733_4_lut_4_lut (.A(n45869), .B(n45923), .C(n45856), 
         .D(n43686), .Z(n45854)) /* synthesis lut_function=(A (B (C+!(D)))+!A !(B ((D)+!C))) */ ;
    defparam i3049_3_lut_rep_733_4_lut_4_lut.init = 16'h91d9;
    LUT4 i24452_4_lut_then_1_lut (.A(akku_o_c_4), .Z(n46335)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i24452_4_lut_then_1_lut.init = 16'h5555;
    LUT4 i24452_4_lut_else_1_lut (.A(akku_o_c_4), .B(akku_o_c_2), .C(akku_o_c_1), 
         .D(akku_o_c_0), .Z(n46334)) /* synthesis lut_function=(!(A (B+(C+(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i24452_4_lut_else_1_lut.init = 16'h5557;
    LUT4 n45315_bdd_3_lut_4_lut_then_4_lut (.A(oprand[2]), .B(oprand[1]), 
         .C(oprand[0]), .D(oprand[4]), .Z(n46338)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+(D)))+!A !(B (C (D))+!B !(C (D)+!C !(D)))) */ ;
    defparam n45315_bdd_3_lut_4_lut_then_4_lut.init = 16'hb66d;
    LUT4 n45315_bdd_3_lut_4_lut_else_4_lut (.A(oprand[2]), .B(oprand[1]), 
         .C(oprand[0]), .D(oprand[4]), .Z(n46337)) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)))+!A (B (C (D)+!C !(D))+!B (C+(D)))) */ ;
    defparam n45315_bdd_3_lut_4_lut_else_4_lut.init = 16'hdbb6;
    LUT4 i2_2_lut_rep_904_4_lut (.A(n46851), .B(n46071), .C(n46850), .D(n46034), 
         .Z(n46025)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_2_lut_rep_904_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_rep_917_3_lut_4_lut_4_lut (.A(n46089), .B(n46078), .C(n130_adj_360), 
         .D(n46091), .Z(n46038)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_rep_917_3_lut_4_lut_4_lut.init = 16'hcdc3;
    LUT4 i37081_4_lut_then_4_lut (.A(n46183), .B(n46264), .C(oprand[3]), 
         .D(oprand[2]), .Z(n46341)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)+!C !(D)))) */ ;
    defparam i37081_4_lut_then_4_lut.init = 16'ha08a;
    CCU2D add_605_5 (.A0(n22564[2]), .B0(n45778), .C0(n46130), .D0(n895[8]), 
          .A1(n45773), .B1(n46130), .C1(n45778), .D1(n895[8]), .CIN(n40505), 
          .COUT(n40506), .S0(n2577[3]), .S1(n2577[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_605_5.INIT0 = 16'h5555;
    defparam add_605_5.INIT1 = 16'h56aa;
    defparam add_605_5.INJECT1_0 = "NO";
    defparam add_605_5.INJECT1_1 = "NO";
    LUT4 i37081_4_lut_else_4_lut (.A(n46183), .B(n46264), .C(oprand[3]), 
         .D(oprand[2]), .Z(n46340)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i37081_4_lut_else_4_lut.init = 16'ha8a0;
    LUT4 i1_4_lut_then_4_lut_adj_94 (.A(oprand[4]), .B(oprand[3]), .C(oprand[0]), 
         .D(oprand[2]), .Z(n46344)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_then_4_lut_adj_94.init = 16'haaa8;
    LUT4 i23730_4_lut (.A(n40788), .B(n46145), .C(n545[0]), .D(n89_adj_320), 
         .Z(n615[0])) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i23730_4_lut.init = 16'h88c0;
    CCU2D add_605_3 (.A0(n43991), .B0(n6_adj_355), .C0(n45778), .D0(GND_net), 
          .A1(n45778), .B1(n46130), .C1(n45776), .D1(n895[8]), .CIN(n40504), 
          .COUT(n40505), .S0(n2577[1]), .S1(n2577[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_605_3.INIT0 = 16'hee1e;
    defparam add_605_3.INIT1 = 16'h6666;
    defparam add_605_3.INJECT1_0 = "NO";
    defparam add_605_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_4_lut (.A(n45898), .B(n41358), .C(n45875), .D(n40960), 
         .Z(n6_adj_361)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_4_lut_4_lut.init = 16'h2bd4;
    LUT4 i37265_2_lut_rep_932_3_lut_4_lut (.A(n46089), .B(n46078), .C(n130_adj_360), 
         .D(n46091), .Z(n46053)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i37265_2_lut_rep_932_3_lut_4_lut.init = 16'hfef0;
    LUT4 i1_4_lut_else_4_lut_adj_95 (.A(oprand[4]), .B(oprand[3]), .C(oprand[2]), 
         .Z(n46343)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i1_4_lut_else_4_lut_adj_95.init = 16'ha8a8;
    LUT4 div_39_i112_3_lut_4_lut_3_lut_4_lut (.A(n46089), .B(n46078), .C(n130_adj_360), 
         .D(n46091), .Z(n161)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_i112_3_lut_4_lut_3_lut_4_lut.init = 16'h11e0;
    LUT4 i37289_3_lut_2_lut_3_lut_4_lut (.A(n46089), .B(n46078), .C(n130_adj_360), 
         .D(n46091), .Z(n160_adj_362)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i37289_3_lut_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 i32417_2_lut_3_lut_4_lut_then_4_lut (.A(oprand[3]), .B(oprand[4]), 
         .C(oprand[2]), .D(oprand[0]), .Z(n46351)) /* synthesis lut_function=(!(A (B (C)+!B !(C+(D)))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam i32417_2_lut_3_lut_4_lut_then_4_lut.init = 16'h3f38;
    LUT4 i32417_2_lut_3_lut_4_lut_else_4_lut (.A(oprand[3]), .B(oprand[4]), 
         .C(oprand[2]), .D(oprand[0]), .Z(n46350)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam i32417_2_lut_3_lut_4_lut_else_4_lut.init = 16'hf8f0;
    LUT4 i38257_then_4_lut (.A(akku_o_c_0), .B(akku_o_c_2), .C(akku_o_c_4), 
         .D(akku_o_c_1), .Z(n46354)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i38257_then_4_lut.init = 16'h2000;
    LUT4 i38257_else_4_lut (.A(akku_o_c_0), .B(akku_o_c_2), .C(akku_o_c_4), 
         .D(akku_o_c_1), .Z(n46353)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i38257_else_4_lut.init = 16'h0001;
    LUT4 div_28_i127_3_lut_4_lut_4_lut (.A(n46088), .B(n12_adj_358), .C(n152), 
         .D(n46073), .Z(n182)) /* synthesis lut_function=(A (C)+!A (B (C (D))+!B (C (D)+!C !(D)))) */ ;
    defparam div_28_i127_3_lut_4_lut_4_lut.init = 16'hf0a1;
    LUT4 div_28_i128_4_lut_rep_937_3_lut_4_lut (.A(n46088), .B(n12_adj_358), 
         .C(n152), .D(n46073), .Z(n46058)) /* synthesis lut_function=(!(A (D)+!A !(B ((D)+!C)+!B (D)))) */ ;
    defparam div_28_i128_4_lut_rep_937_3_lut_4_lut.init = 16'h55ae;
    LUT4 i1_4_lut_3_lut_4_lut_then_4_lut (.A(akku_o_c_4), .B(akku_o_c_1), 
         .C(akku_o_c_2), .D(akku_o_c_3), .Z(n46357)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i1_4_lut_3_lut_4_lut_then_4_lut.init = 16'h1400;
    LUT4 i1_4_lut_3_lut_4_lut_else_4_lut (.A(akku_o_c_4), .B(akku_o_c_2), 
         .C(akku_o_c_3), .Z(n46356)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i1_4_lut_3_lut_4_lut_else_4_lut.init = 16'h4040;
    LUT4 div_39_i113_3_lut_rep_918_4_lut_4_lut (.A(n46089), .B(n46078), 
         .C(n46091), .D(n130_adj_360), .Z(n46039)) /* synthesis lut_function=(A (B+!(C+(D)))+!A !(B+!(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_i113_3_lut_rep_918_4_lut_4_lut.init = 16'h998a;
    LUT4 mux_47_i6_3_lut_rep_913_4_lut (.A(n46079), .B(n46093), .C(n46123), 
         .D(n46042), .Z(n46034)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_47_i6_3_lut_rep_913_4_lut.init = 16'hfe0e;
    LUT4 i4988_4_lut_then_4_lut (.A(n2203[5]), .B(n45757), .C(n43670), 
         .D(n790[4]), .Z(n46360)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i4988_4_lut_then_4_lut.init = 16'h19da;
    LUT4 i4988_4_lut_else_4_lut (.A(n2203[5]), .B(n45757), .C(n43670), 
         .D(n790[4]), .Z(n46359)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A (B ((D)+!C)+!B !(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i4988_4_lut_else_4_lut.init = 16'h185a;
    LUT4 i2_3_lut_4_lut_adj_96 (.A(n45874), .B(n45921), .C(n22874), .D(n45865), 
         .Z(n23447)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_4_lut_adj_96.init = 16'h0f78;
    LUT4 i15159_3_lut_rep_633 (.A(n790[4]), .B(n2203[5]), .C(n45757), 
         .Z(n45754)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i15159_3_lut_rep_633.init = 16'ha8a8;
    LUT4 i4953_4_lut_then_4_lut (.A(n45762), .B(n2203[5]), .C(n2072[5]), 
         .D(n790[4]), .Z(n46363)) /* synthesis lut_function=(A (B (D))+!A (B+!(C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i4953_4_lut_then_4_lut.init = 16'hcd44;
    LUT4 i4953_4_lut_else_4_lut (.A(n45762), .B(n2203[5]), .C(n755[3]), 
         .D(n790[4]), .Z(n46362)) /* synthesis lut_function=(A (B (D))+!A (B+(C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i4953_4_lut_else_4_lut.init = 16'hdc44;
    LUT4 div_28_i126_4_lut_4_lut (.A(n46088), .B(n12_adj_358), .C(n152), 
         .D(n46065), .Z(n181)) /* synthesis lut_function=(!(A (C+(D))+!A (B+(C+(D))))) */ ;
    defparam div_28_i126_4_lut_4_lut.init = 16'h000b;
    LUT4 i34_4_lut_4_lut_then_4_lut (.A(n46160), .B(akku_o_c_2), .C(akku_o_c_3), 
         .D(akku_o_c_4), .Z(n46366)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C+(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i34_4_lut_4_lut_then_4_lut.init = 16'h5154;
    LUT4 i34_4_lut_4_lut_else_4_lut (.A(n46160), .B(akku_o_c_2), .C(akku_o_c_3), 
         .D(akku_o_c_4), .Z(n46365)) /* synthesis lut_function=(!(A+!(B (C)+!B !(C (D)+!C !(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i34_4_lut_4_lut_else_4_lut.init = 16'h4150;
    LUT4 i38254_then_3_lut (.A(oprand[2]), .B(oprand[3]), .C(oprand[1]), 
         .Z(n46369)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i38254_then_3_lut.init = 16'h0101;
    LUT4 i23729_4_lut (.A(n46400), .B(n46128), .C(n475[0]), .D(n45_adj_356), 
         .Z(n545[0])) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i23729_4_lut.init = 16'h88c0;
    LUT4 i38254_else_3_lut (.A(oprand[2]), .B(oprand[3]), .C(oprand[0]), 
         .D(oprand[1]), .Z(n46368)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i38254_else_3_lut.init = 16'h0001;
    LUT4 mux_160_i4_3_lut_rep_1161 (.A(n1829[5]), .B(n685[3]), .C(n89), 
         .Z(n46847)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_160_i4_3_lut_rep_1161.init = 16'h5c5c;
    LUT4 i2_4_lut_then_4_lut_adj_97 (.A(n45823), .B(n46051), .C(n45885), 
         .D(n45794), .Z(n46372)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(C+(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_4_lut_then_4_lut_adj_97.init = 16'h3336;
    LUT4 i2_4_lut_else_4_lut (.A(n45823), .B(n89_adj_303), .C(n45829), 
         .D(n45885), .Z(n46371)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (B+((D)+!C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_4_lut_else_4_lut.init = 16'hff65;
    LUT4 i14941_3_lut_4_lut (.A(n45874), .B(n45921), .C(n45865), .D(n22874), 
         .Z(n4_adj_363)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i14941_3_lut_4_lut.init = 16'h00f8;
    LUT4 i38246_then_4_lut (.A(oprand[4]), .B(oprand[3]), .C(oprand[0]), 
         .D(oprand[1]), .Z(n46375)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i38246_then_4_lut.init = 16'h0020;
    LUT4 i38234_then_4_lut (.A(akku_o_c_3), .B(akku_o_c_2), .C(akku_o_c_0), 
         .D(akku_o_c_1), .Z(n46378)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(C+(D))))) */ ;
    defparam i38234_then_4_lut.init = 16'h4001;
    LUT4 i1_3_lut_rep_943_4_lut (.A(n46084), .B(n46096), .C(n29_adj_353), 
         .D(n46851), .Z(n46064)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_3_lut_rep_943_4_lut.init = 16'h8f00;
    LUT4 i1_2_lut_rep_630_4_lut (.A(n790[4]), .B(n2203[5]), .C(n45757), 
         .D(n45762), .Z(n45751)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_rep_630_4_lut.init = 16'h57a8;
    LUT4 i1_4_lut_then_4_lut_adj_98 (.A(n18[5]), .B(n18[3]), .C(n18[2]), 
         .D(n257), .Z(n46381)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;
    defparam i1_4_lut_then_4_lut_adj_98.init = 16'heeea;
    LUT4 i1_4_lut_else_4_lut_adj_99 (.A(n45974), .B(n45981), .C(n45982), 
         .D(n257), .Z(n46380)) /* synthesis lut_function=(A (B+!(C))+!A (B+!(C+!(D)))) */ ;
    defparam i1_4_lut_else_4_lut_adj_99.init = 16'hcfce;
    LUT4 i3_4_lut_rep_1167 (.A(data[5]), .B(akku_o_c_8), .C(data[6]), 
         .D(data[7]), .Z(n46853)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i3_4_lut_rep_1167.init = 16'h4000;
    LUT4 i2_4_lut_adj_100 (.A(n21411), .B(n46036), .C(n6324), .D(n4_adj_317), 
         .Z(n22855)) /* synthesis lut_function=(A (B+(D))+!A (B (C)+!B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_4_lut_adj_100.init = 16'hfac9;
    LUT4 i38232_then_4_lut (.A(oprand[4]), .B(oprand[3]), .C(oprand[0]), 
         .D(oprand[1]), .Z(n46384)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i38232_then_4_lut.init = 16'h2000;
    LUT4 i38232_else_4_lut (.A(oprand[3]), .B(oprand[0]), .C(oprand[1]), 
         .Z(n46383)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i38232_else_4_lut.init = 16'h0101;
    LUT4 n45395_bdd_3_lut_then_4_lut (.A(oprand[0]), .B(oprand[3]), .C(oprand[2]), 
         .D(akku_o_c_2), .Z(n46387)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam n45395_bdd_3_lut_then_4_lut.init = 16'h0008;
    LUT4 n45395_bdd_3_lut_else_4_lut (.A(oprand[0]), .B(oprand[3]), .C(oprand[2]), 
         .D(akku_o_c_2), .Z(n46386)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam n45395_bdd_3_lut_else_4_lut.init = 16'h0800;
    LUT4 i5486_3_lut_3_lut_rep_608_4_lut (.A(n44713), .B(n45732), .C(n45735), 
         .D(n45728), .Z(n45729)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5486_3_lut_3_lut_rep_608_4_lut.init = 16'hf069;
    LUT4 n107_bdd_4_lut_then_4_lut (.A(oprand[0]), .B(oprand[2]), .C(oprand[3]), 
         .D(oprand[1]), .Z(n46390)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (((D)+!C)+!B))) */ ;
    defparam n107_bdd_4_lut_then_4_lut.init = 16'h0048;
    LUT4 i1_4_lut_4_lut (.A(akku_o_c_4), .B(akku_o_c_3), .C(akku_o_c_2), 
         .D(akku_o_c_1), .Z(n9)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i1_4_lut_4_lut.init = 16'h0002;
    CCU2D add_275_5 (.A0(n475[8]), .B0(n46035), .C0(n38153), .D0(n23007), 
          .A1(n43902), .B1(n46035), .C1(n30789), .D1(n16[8]), .CIN(n40420), 
          .COUT(n40421), .S0(n999[3]), .S1(n999[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_275_5.INIT0 = 16'hf00f;
    defparam add_275_5.INIT1 = 16'h5555;
    defparam add_275_5.INJECT1_0 = "NO";
    defparam add_275_5.INJECT1_1 = "NO";
    LUT4 n107_bdd_4_lut_else_4_lut (.A(oprand[0]), .B(oprand[2]), .C(oprand[3]), 
         .D(oprand[1]), .Z(n46389)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C (D))+!B !(C+(D))))) */ ;
    defparam n107_bdd_4_lut_else_4_lut.init = 16'h4801;
    LUT4 n100_bdd_4_lut_4_lut (.A(n46096), .B(n46083), .C(n46123), .D(n46097), 
         .Z(n130)) /* synthesis lut_function=(!((B ((D)+!C)+!B !(C))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam n100_bdd_4_lut_4_lut.init = 16'h20a0;
    LUT4 akku_o_c_0_bdd_4_lut_38209 (.A(akku_o_c_0), .B(n46271), .C(n46248), 
         .D(akku_o_c_1), .Z(n31204)) /* synthesis lut_function=(A (B (C+!(D))+!B (C+(D)))+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam akku_o_c_0_bdd_4_lut_38209.init = 16'hf2ec;
    LUT4 i23724_2_lut_rep_1171 (.A(n46882), .B(n46880), .Z(n46870)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23724_2_lut_rep_1171.init = 16'heeee;
    LUT4 n45474_bdd_2_lut (.A(n45474), .B(n930[1]), .Z(n45475)) /* synthesis lut_function=(A+(B)) */ ;
    defparam n45474_bdd_2_lut.init = 16'heeee;
    LUT4 i23900_2_lut_3_lut_4_lut (.A(data[5]), .B(akku_o_c_8), .C(data[6]), 
         .D(data[7]), .Z(states_2__N_76[2])) /* synthesis lut_function=(A (D)+!A (B (C (D)))) */ ;
    defparam i23900_2_lut_3_lut_4_lut.init = 16'hea00;
    FD1S3IX states__i2 (.D(states_2__N_76[2]), .CK(clk_c), .CD(n46244), 
            .Q(states_c[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam states__i2.GSR = "ENABLED";
    FD1S3AX adreg_i1 (.D(adress_5__N_3[1]), .CK(clk_c), .Q(address[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam adreg_i1.GSR = "ENABLED";
    LUT4 i5570_3_lut (.A(n2629[0]), .B(n2629[5]), .C(n895[0]), .Z(n2_adj_367)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5570_3_lut.init = 16'hb2b2;
    LUT4 i1_4_lut_then_4_lut_adj_101 (.A(n108_adj_368), .B(n270[5]), .C(n270[2]), 
         .D(n270[1]), .Z(n46396)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i1_4_lut_then_4_lut_adj_101.init = 16'heccc;
    LUT4 i1_4_lut_else_4_lut_adj_102 (.A(n108_adj_368), .B(n253), .C(n107_adj_346), 
         .D(n256), .Z(n46395)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i1_4_lut_else_4_lut_adj_102.init = 16'heccc;
    LUT4 n1147_bdd_4_lut_38317 (.A(n45896), .B(n46051), .C(n45829), .D(n46122), 
         .Z(n6_adj_369)) /* synthesis lut_function=(A (B+!(D))+!A ((C+!(D))+!B)) */ ;
    defparam n1147_bdd_4_lut_38317.init = 16'hd9ff;
    LUT4 i2_3_lut_4_lut_4_lut_4_lut (.A(n45779), .B(n860[5]), .C(n45758), 
         .D(n45743), .Z(n2476[3])) /* synthesis lut_function=(A (B (C)+!B !(C (D)))+!A (B (C (D))+!B !(C (D)))) */ ;
    defparam i2_3_lut_4_lut_4_lut_4_lut.init = 16'hc3b3;
    LUT4 i2_4_lut_then_4_lut_adj_103 (.A(n1051[5]), .B(n1051[4]), .C(n1051[2]), 
         .D(n4_adj_370), .Z(n46399)) /* synthesis lut_function=(A (B)+!A !(B (C+(D))+!B !(C+(D)))) */ ;
    defparam i2_4_lut_then_4_lut_adj_103.init = 16'h999c;
    LUT4 i2_4_lut_else_4_lut_adj_104 (.A(n1051[5]), .B(n1051[4]), .C(n1051[2]), 
         .D(n4_adj_370), .Z(n46398)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A (B)) */ ;
    defparam i2_4_lut_else_4_lut_adj_104.init = 16'hc666;
    LUT4 mux_107_i1_4_lut (.A(n7_adj_371), .B(n429[0]), .C(n37), .D(n8_adj_372), 
         .Z(n462[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !(B (C (D))+!B ((D)+!C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_107_i1_4_lut.init = 16'hac5c;
    LUT4 i2_4_lut_adj_105 (.A(n41383), .B(n6_adj_373), .C(n9938), .D(n21933), 
         .Z(n7_adj_371)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C+(D))+!B !(C+(D))))) */ ;
    defparam i2_4_lut_adj_105.init = 16'h393c;
    LUT4 i38137_4_lut (.A(akku_o_c_4), .B(n43941), .C(n77), .D(n46223), 
         .Z(n44765)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B+!(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i38137_4_lut.init = 16'hcfef;
    LUT4 i24472_4_lut_then_4_lut (.A(oprand[4]), .B(oprand[3]), .C(oprand[2]), 
         .D(oprand[1]), .Z(n46402)) /* synthesis lut_function=(!(A (B+(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam i24472_4_lut_then_4_lut.init = 16'h5777;
    PFUMX i38437 (.BLUT(n46293), .ALUT(n46294), .C0(n46205), .Z(n51_adj_345));
    LUT4 mux_195_i6_3_lut_4_lut (.A(n45779), .B(n860[5]), .C(n45758), 
         .D(n46157), .Z(n895[5])) /* synthesis lut_function=(A (B (C+(D)))+!A (B (D))) */ ;
    defparam mux_195_i6_3_lut_4_lut.init = 16'hcc80;
    LUT4 i2_4_lut_then_4_lut_adj_106 (.A(akku_o_c_0), .B(akku_o_c_4), .C(akku_o_c_2), 
         .D(akku_o_c_3), .Z(n46858)) /* synthesis lut_function=(!((B (C+!(D))+!B !(C))+!A)) */ ;
    defparam i2_4_lut_then_4_lut_adj_106.init = 16'h2820;
    LUT4 i2_4_lut_then_4_lut_adj_107 (.A(n1582[5]), .B(n1582[4]), .C(n1582[2]), 
         .D(n4_adj_374), .Z(n46405)) /* synthesis lut_function=(A (B)+!A !(B (C+(D))+!B !(C+(D)))) */ ;
    defparam i2_4_lut_then_4_lut_adj_107.init = 16'h999c;
    LUT4 i1_2_lut_3_lut_4_lut_adj_108 (.A(n45877), .B(n45920), .C(n43689), 
         .D(n45921), .Z(n541[4])) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (C)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_3_lut_4_lut_adj_108.init = 16'hd2f0;
    LUT4 i2_4_lut_else_4_lut_adj_109 (.A(n1582[5]), .B(n1582[4]), .C(n1582[2]), 
         .D(n4_adj_374), .Z(n46404)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A (B)) */ ;
    defparam i2_4_lut_else_4_lut_adj_109.init = 16'hc666;
    LUT4 i63_then_4_lut (.A(akku_o_c_0), .B(n46191), .C(n117_adj_305), 
         .D(n122_adj_375), .Z(n46288)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i63_then_4_lut.init = 16'h2000;
    LUT4 i1_3_lut_4_lut_adj_110 (.A(n45779), .B(n860[5]), .C(n45758), 
         .D(n45743), .Z(n2476[2])) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_110.init = 16'h0f70;
    LUT4 mux_174_i4_3_lut_rep_636 (.A(n2072[5]), .B(n755[3]), .C(n43564), 
         .Z(n45757)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_174_i4_3_lut_rep_636.init = 16'h5c5c;
    LUT4 i2589_4_lut_then_4_lut (.A(n405[2]), .B(n45929), .C(n45940), 
         .D(n293[1]), .Z(n46408)) /* synthesis lut_function=(A (B+!(D))+!A !((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2589_4_lut_then_4_lut.init = 16'h8cae;
    CCU2D add_275_3 (.A0(n45900), .B0(n475[8]), .C0(n46035), .D0(n46017), 
          .A1(n45900), .B1(n46035), .C1(n475[8]), .D1(n46017), .CIN(n40419), 
          .COUT(n40420), .S0(n999[1]), .S1(n999[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_275_3.INIT0 = 16'ha956;
    defparam add_275_3.INIT1 = 16'h659a;
    defparam add_275_3.INJECT1_0 = "NO";
    defparam add_275_3.INJECT1_1 = "NO";
    LUT4 i63_else_4_lut (.A(akku_o_c_0), .B(n46191), .C(n117_adj_305), 
         .D(n122_adj_375), .Z(n46287)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i63_else_4_lut.init = 16'h0001;
    LUT4 i2589_4_lut_else_4_lut (.A(n405[2]), .B(n45929), .C(n3[4]), .D(n45940), 
         .Z(n46407)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2589_4_lut_else_4_lut.init = 16'heaa8;
    CCU2D add_605_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n45758), .B1(n45779), .C1(n46157), .D1(n860[5]), .COUT(n40504), 
          .S1(n2577[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_605_1.INIT0 = 16'hF000;
    defparam add_605_1.INIT1 = 16'h07ff;
    defparam add_605_1.INJECT1_0 = "NO";
    defparam add_605_1.INJECT1_1 = "NO";
    LUT4 n1688_bdd_4_lut (.A(n1687[5]), .B(n45794), .C(n45823), .D(n45790), 
         .Z(n6_adj_376)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A !(B+(C))) */ ;
    defparam n1688_bdd_4_lut.init = 16'ha383;
    LUT4 i2311_4_lut_3_lut_rep_754 (.A(n41358), .B(n45902), .C(n45909), 
         .Z(n45875)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2311_4_lut_3_lut_rep_754.init = 16'h8e8e;
    LUT4 i23728_4_lut (.A(n43766), .B(n15_adj_316), .C(n363[0]), .D(n37_adj_301), 
         .Z(n429[0])) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C+(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i23728_4_lut.init = 16'h44c0;
    LUT4 i4_4_lut (.A(n41360), .B(n43765), .C(n45824), .D(n6_adj_377), 
         .Z(n43766)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i4_4_lut.init = 16'h6996;
    LUT4 i1_4_lut_adj_111 (.A(n22740), .B(n6_adj_378), .C(n9966), .D(n21939), 
         .Z(n6_adj_377)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A (B (C)+!B !(C)))) */ ;
    defparam i1_4_lut_adj_111.init = 16'h363c;
    LUT4 i1_2_lut_rep_632_4_lut (.A(n2072[5]), .B(n755[3]), .C(n43564), 
         .D(n2203[5]), .Z(n45753)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(B (D)+!B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_632_4_lut.init = 16'ha35c;
    LUT4 i2_3_lut_rep_945_4_lut (.A(n46086), .B(n46196), .C(n45_adj_356), 
         .D(n46128), .Z(n46066)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i2_3_lut_rep_945_4_lut.init = 16'h0800;
    LUT4 i5850_4_lut (.A(n45842), .B(n9959), .C(n21937), .D(n4_adj_379), 
         .Z(n4_adj_380)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B+(C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5850_4_lut.init = 16'hdcec;
    LUT4 n587_bdd_4_lut (.A(n580[2]), .B(n580[1]), .C(n1429[1]), .D(n45796), 
         .Z(n45547)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;
    defparam n587_bdd_4_lut.init = 16'h5e8f;
    LUT4 i23727_4_lut (.A(n43769), .B(n15), .C(n3[0]), .D(n37_adj_340), 
         .Z(n363[0])) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i23727_4_lut.init = 16'h88c0;
    LUT4 i6_4_lut (.A(n11_adj_381), .B(n9_adj_382), .C(n22902), .D(n45870), 
         .Z(n43769)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i6_4_lut.init = 16'h6996;
    LUT4 i4_3_lut (.A(n43768), .B(n41385), .C(n41077), .Z(n11_adj_381)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;
    defparam i4_3_lut.init = 16'h6969;
    LUT4 i2_4_lut_adj_112 (.A(n6_adj_321), .B(n40744), .C(n42171), .D(n44079), 
         .Z(n9_adj_382)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A !(B (C)+!B (C+(D))))) */ ;
    defparam i2_4_lut_adj_112.init = 16'h595a;
    LUT4 i23859_2_lut_rep_938_3_lut_4_lut (.A(n37_adj_301), .B(n46087), 
         .C(n46136), .D(n15_adj_316), .Z(n46059)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i23859_2_lut_rep_938_3_lut_4_lut.init = 16'h4000;
    LUT4 i17142_2_lut_rep_939_3_lut_4_lut (.A(n37_adj_301), .B(n46087), 
         .C(n37), .D(n15_adj_316), .Z(n46060)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i17142_2_lut_rep_939_3_lut_4_lut.init = 16'h0400;
    LUT4 i2_3_lut (.A(n3[1]), .B(n41242), .C(n3[2]), .Z(n41411)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i2_3_lut.init = 16'h9696;
    LUT4 i1_2_lut_rep_749_4_lut_4_lut (.A(n3[4]), .B(n45880), .C(n3[3]), 
         .D(n22900), .Z(n45870)) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_rep_749_4_lut_4_lut.init = 16'h8e71;
    LUT4 i23726_4_lut (.A(n41374), .B(n43592), .C(n231_adj_515[0]), .D(n37_adj_318), 
         .Z(n3[0])) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B+!(C+(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i23726_4_lut.init = 16'h1130;
    LUT4 i4_4_lut_adj_113 (.A(n41358), .B(n6_adj_383), .C(n41402), .D(n6_adj_361), 
         .Z(n41374)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i4_4_lut_adj_113.init = 16'h9669;
    LUT4 i5913_4_lut (.A(n45875), .B(n10022), .C(n21951), .D(n4_adj_384), 
         .Z(n6_adj_383)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B+(C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5913_4_lut.init = 16'hdcec;
    LUT4 i1_4_lut_adj_114 (.A(n43581), .B(n46048), .C(n22585), .D(n46104), 
         .Z(n825[7])) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_114.init = 16'h8000;
    LUT4 i3013_2_lut_3_lut_3_lut_rep_797_4_lut (.A(n46136), .B(n46087), 
         .C(n45869), .D(n45923), .Z(n45918)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(D)) */ ;
    defparam i3013_2_lut_3_lut_3_lut_rep_797_4_lut.init = 16'h88f7;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(n46136), .B(n46087), .C(n45869), 
         .D(n45923), .Z(n43675)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'h7778;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n3[4]), .B(n45880), .C(n3[3]), 
         .D(n22900), .Z(n22894)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h42bd;
    LUT4 i2_3_lut_rep_920_4_lut (.A(n89_adj_303), .B(n46055), .C(n46137), 
         .D(n43547), .Z(n46041)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i2_3_lut_rep_920_4_lut.init = 16'h4000;
    LUT4 i14923_3_lut_rep_750_4_lut_4_lut (.A(n3[4]), .B(n45880), .C(n3[3]), 
         .D(n22900), .Z(n45871)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i14923_3_lut_rep_750_4_lut_4_lut.init = 16'h00fd;
    LUT4 i2623_2_lut_3_lut_4_lut_4_lut (.A(n3[4]), .B(n45880), .C(n3[3]), 
         .D(n22900), .Z(n6734)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2623_2_lut_3_lut_4_lut_4_lut.init = 16'h0031;
    LUT4 akku_o_c_4_bdd_4_lut_38441 (.A(akku_o_c_4), .B(akku_o_c_3), .C(akku_o_c_2), 
         .D(akku_o_c_1), .Z(n9_adj_385)) /* synthesis lut_function=(!((B (C (D)))+!A)) */ ;
    defparam akku_o_c_4_bdd_4_lut_38441.init = 16'h2aaa;
    LUT4 i1_2_lut_adj_115 (.A(n45287), .B(n45286), .Z(n29_adj_353)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_2_lut_adj_115.init = 16'h8888;
    LUT4 i5155_2_lut_rep_631_4_lut (.A(n2332[5]), .B(n825[4]), .C(n45), 
         .D(n860[5]), .Z(n45752)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(B (D)+!B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i5155_2_lut_rep_631_4_lut.init = 16'ha35c;
    LUT4 i2775_2_lut_rep_753_4_lut (.A(n45880), .B(n3[4]), .C(n37_adj_340), 
         .D(n45920), .Z(n45874)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A ((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i2775_2_lut_rep_753_4_lut.init = 16'h00ac;
    LUT4 i1_2_lut_4_lut_adj_116 (.A(n45880), .B(n3[4]), .C(n37_adj_340), 
         .D(n45920), .Z(n22874)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_4_lut_adj_116.init = 16'h53ac;
    LUT4 i5160_2_lut_4_lut (.A(n2332[5]), .B(n825[4]), .C(n45), .D(n860[5]), 
         .Z(n4_adj_386)) /* synthesis lut_function=(!(A (B (C (D))+!B (D))+!A !(B+(C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i5160_2_lut_4_lut.init = 16'h5cff;
    LUT4 i2_4_lut_4_lut_adj_117 (.A(n1855[3]), .B(n1855[5]), .C(n6_adj_350), 
         .D(n1855[4]), .Z(n40781)) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_4_lut_4_lut_adj_117.init = 16'hdb24;
    LUT4 i1_2_lut_rep_602_4_lut (.A(n2616[5]), .B(n895[2]), .C(n43563), 
         .D(n45727), .Z(n45723)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A (B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_602_4_lut.init = 16'hff5c;
    LUT4 mux_167_i5_3_lut_4_lut (.A(n45765), .B(n45760), .C(n19), .D(n45791), 
         .Z(n755[4])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_167_i5_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_58_i1_3_lut (.A(n218[3]), .B(n218[0]), .C(n46179), .Z(n231_adj_515[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_58_i1_3_lut.init = 16'hcaca;
    CCU2D add_559_7 (.A0(n2358[4]), .B0(n2358[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40503), 
          .S0(n2371[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_559_7.INIT0 = 16'h5999;
    defparam add_559_7.INIT1 = 16'h0000;
    defparam add_559_7.INJECT1_0 = "NO";
    defparam add_559_7.INJECT1_1 = "NO";
    LUT4 i6463_2_lut_rep_909_3_lut_4_lut (.A(n46069), .B(n130_adj_360), 
         .C(n46050), .D(n46078), .Z(n46030)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C+(D)))) */ ;
    defparam i6463_2_lut_rep_909_3_lut_4_lut.init = 16'hf1fe;
    LUT4 mux_54_i1_4_lut (.A(n11_adj_388), .B(n108_adj_368), .C(n29_adj_353), 
         .D(n45663), .Z(n218[0])) /* synthesis lut_function=(A (B+(C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_54_i1_4_lut.init = 16'hfcac;
    LUT4 i4_4_lut_adj_118 (.A(n45912), .B(n46397), .C(n270[6]), .D(n208[1]), 
         .Z(n11_adj_388)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;
    defparam i4_4_lut_adj_118.init = 16'hfcee;
    LUT4 i5675_4_lut_3_lut (.A(n1855[5]), .B(n685[0]), .C(n1855[0]), .Z(n2_adj_349)) /* synthesis lut_function=(A (B+(C))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5675_4_lut_3_lut.init = 16'he8e8;
    LUT4 i1_2_lut_rep_931_4_lut (.A(n46145), .B(n89_adj_320), .C(n46066), 
         .D(n89_adj_303), .Z(n46052)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_931_4_lut.init = 16'h0020;
    LUT4 i4692_4_lut_rep_640 (.A(n1947[2]), .B(n45764), .C(n23877), .D(n45770), 
         .Z(n45761)) /* synthesis lut_function=(A (B+(C))+!A !((D)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i4692_4_lut_rep_640.init = 16'ha8ec;
    LUT4 i6554_2_lut_rep_910_4_lut_4_lut_4_lut (.A(n46092), .B(n46083), 
         .C(n46093), .D(n46042), .Z(n46031)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))+!B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i6554_2_lut_rep_910_4_lut_4_lut_4_lut.init = 16'h7662;
    LUT4 i4697_2_lut_rep_639_3_lut (.A(n1947[2]), .B(n45764), .C(n45770), 
         .Z(n45760)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i4697_2_lut_rep_639_3_lut.init = 16'h8c8c;
    LUT4 i14976_3_lut_4_lut (.A(n23650), .B(n46082), .C(n46019), .D(n43592), 
         .Z(n4201[1])) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((D)+!C))) */ ;
    defparam i14976_3_lut_4_lut.init = 16'h0078;
    LUT4 i1_2_lut_4_lut_4_lut_adj_119 (.A(n45881), .B(n4217[1]), .C(n45883), 
         .D(n4_adj_389), .Z(n40857)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_119.init = 16'h5955;
    LUT4 i24246_2_lut_3_lut_4_lut (.A(n23650), .B(n46082), .C(n43592), 
         .D(n46019), .Z(n6383)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i24246_2_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 i14924_3_lut_rep_755_4_lut (.A(n45929), .B(n43720), .C(n3[3]), 
         .D(n3[4]), .Z(n45876)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A (B ((D)+!C)+!B (D)))) */ ;
    defparam i14924_3_lut_rep_755_4_lut.init = 16'h00f9;
    LUT4 mux_174_i6_3_lut_rep_641 (.A(n2046[5]), .B(n755[5]), .C(n43564), 
         .Z(n45762)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_174_i6_3_lut_rep_641.init = 16'h5c5c;
    LUT4 mux_79_i5_3_lut_rep_756_4_lut (.A(n45929), .B(n43720), .C(n37_adj_340), 
         .D(n3[4]), .Z(n45877)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_79_i5_3_lut_rep_756_4_lut.init = 16'h6f60;
    CCU2D add_559_5 (.A0(n2358[2]), .B0(n2358[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2358[3]), .B1(n2358[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40502), .COUT(n40503), .S0(n2371[3]), .S1(n2371[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_559_5.INIT0 = 16'h5666;
    defparam add_559_5.INIT1 = 16'h5666;
    defparam add_559_5.INJECT1_0 = "NO";
    defparam add_559_5.INJECT1_1 = "NO";
    LUT4 mux_195_i3_4_lut_4_lut (.A(n45731), .B(n43712), .C(n46157), .D(n45738), 
         .Z(n895[2])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_195_i3_4_lut_4_lut.init = 16'hf606;
    LUT4 i5605_4_lut_3_lut (.A(n2371[5]), .B(n825[0]), .C(n2371[0]), .Z(n2_adj_390)) /* synthesis lut_function=(A (B+(C))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5605_4_lut_3_lut.init = 16'he8e8;
    LUT4 mux_47_i1_4_lut (.A(n30878), .B(n108), .C(n46123), .D(n43333), 
         .Z(n108_adj_368)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_47_i1_4_lut.init = 16'hcfca;
    LUT4 mux_58_i5_3_lut_rep_826_4_lut (.A(n46136), .B(n46095), .C(n46179), 
         .D(n218[4]), .Z(n45947)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam mux_58_i5_3_lut_rep_826_4_lut.init = 16'hf808;
    LUT4 i2_3_lut_4_lut_adj_120 (.A(n45929), .B(n43720), .C(n3[4]), .D(n3[3]), 
         .Z(n427[1])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i2_3_lut_4_lut_adj_120.init = 16'h6996;
    LUT4 mux_160_i3_3_lut_rep_642 (.A(n1842[5]), .B(n685[2]), .C(n89), 
         .Z(n45763)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_160_i3_3_lut_rep_642.init = 16'h5c5c;
    LUT4 mux_188_i6_4_lut (.A(n2319[5]), .B(n45762), .C(n45), .D(n46138), 
         .Z(n860[5])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C+(D))+!B (C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_188_i6_4_lut.init = 16'h5c50;
    CCU2D add_559_3 (.A0(n2358[0]), .B0(n2358[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2358[1]), .B1(n2358[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40501), .COUT(n40502), .S0(n2371[1]), .S1(n2371[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_559_3.INIT0 = 16'h5666;
    defparam add_559_3.INIT1 = 16'h5999;
    defparam add_559_3.INJECT1_0 = "NO";
    defparam add_559_3.INJECT1_1 = "NO";
    LUT4 i17131_2_lut_4_lut (.A(n1842[5]), .B(n685[2]), .C(n89), .D(n45770), 
         .Z(n23877)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B (D)+!B ((D)+!C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i17131_2_lut_4_lut.init = 16'h005c;
    CCU2D add_559_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n43710), .B1(n7_adj_392), .C1(n46138), .D1(n790[1]), .COUT(n40501), 
          .S1(n2371[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_559_1.INIT0 = 16'hF000;
    defparam add_559_1.INIT1 = 16'h09f9;
    defparam add_559_1.INJECT1_0 = "NO";
    defparam add_559_1.INJECT1_1 = "NO";
    LUT4 i23755_3_lut_4_lut (.A(n46136), .B(n46095), .C(n46179), .D(n46090), 
         .Z(n4_adj_317)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i23755_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_153_i2_4_lut_4_lut (.A(n45766), .B(n46137), .C(n650[1]), 
         .D(n40913), .Z(n685[1])) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (B (C)+!B (D))) */ ;
    defparam mux_153_i2_4_lut_4_lut.init = 16'hd1e2;
    LUT4 n6_bdd_3_lut_4_lut (.A(n45789), .B(n45787), .C(n1947[2]), .D(n45763), 
         .Z(n45633)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam n6_bdd_3_lut_4_lut.init = 16'h87f0;
    LUT4 i1_2_lut_adj_121 (.A(n19), .B(n89), .Z(n43547)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_adj_121.init = 16'h2222;
    LUT4 i1_3_lut_4_lut_4_lut_adj_122 (.A(n45908), .B(n46848), .C(n21[2]), 
         .D(n43759), .Z(n4_adj_393)) /* synthesis lut_function=(A (B (C (D))+!B !(C+(D)))+!A !(B (C+!(D))+!B ((D)+!C))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_122.init = 16'h8412;
    LUT4 mux_72_i4_3_lut_4_lut (.A(n45908), .B(n46848), .C(n43592), .D(n45899), 
         .Z(n3[3])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_72_i4_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_174_i5_3_lut (.A(n2059[5]), .B(n755[4]), .C(n43564), .Z(n790[4])) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_174_i5_3_lut.init = 16'h5c5c;
    LUT4 i4854_2_lut_4_lut (.A(n46090), .B(n46041), .C(n43581), .D(n825[7]), 
         .Z(n8965)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i4854_2_lut_4_lut.init = 16'h8000;
    LUT4 n305_bdd_4_lut_4_lut (.A(n45908), .B(n46848), .C(n45899), .D(n45910), 
         .Z(n45583)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;
    defparam n305_bdd_4_lut_4_lut.init = 16'h05e2;
    LUT4 i6938_2_lut_rep_958_4_lut (.A(n46101), .B(n102), .C(n11), .D(n46092), 
         .Z(n46079)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i6938_2_lut_rep_958_4_lut.init = 16'hca00;
    LUT4 i2_3_lut_rep_719_4_lut (.A(n545[8]), .B(n45886), .C(n4217[1]), 
         .D(n4_adj_389), .Z(n45840)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+!(C (D)))) */ ;
    defparam i2_3_lut_rep_719_4_lut.init = 16'h9000;
    LUT4 n41077_bdd_4_lut (.A(n41242), .B(n45851), .C(n45858), .D(n45853), 
         .Z(n45568)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(C)) */ ;
    defparam n41077_bdd_4_lut.init = 16'ha587;
    LUT4 i2_2_lut_4_lut_4_lut (.A(oprand[3]), .B(n46878), .C(oprand[2]), 
         .D(oprand[4]), .Z(n8_adj_394)) /* synthesis lut_function=(A (B+(C+!(D)))+!A !(B+(C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam i2_2_lut_4_lut_4_lut.init = 16'ha9aa;
    LUT4 i31576_2_lut_rep_697_3_lut_4_lut_3_lut_4_lut (.A(n4382[1]), .B(n45884), 
         .C(n38297), .D(n4382[2]), .Z(n45818)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B !(C+(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i31576_2_lut_rep_697_3_lut_4_lut_3_lut_4_lut.init = 16'h1ffe;
    LUT4 i31573_2_lut_rep_699_3_lut_4_lut (.A(n4382[1]), .B(n45884), .C(n38297), 
         .D(n4382[2]), .Z(n45820)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i31573_2_lut_rep_699_3_lut_4_lut.init = 16'hf1fe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_123 (.A(n46098), .B(n37), .C(n46090), 
         .D(n46196), .Z(n475[8])) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_3_lut_4_lut_adj_123.init = 16'h2000;
    LUT4 i1_2_lut_4_lut_4_lut_adj_124 (.A(n45887), .B(n45888), .C(n1403[1]), 
         .D(n46145), .Z(n40970)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A !(B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_124.init = 16'ha595;
    LUT4 i24062_2_lut_3_lut_4_lut (.A(n46098), .B(n37), .C(n46100), .D(n46196), 
         .Z(n30789)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i24062_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 n728_bdd_3_lut_4_lut (.A(n45789), .B(n45787), .C(n45770), .D(n45763), 
         .Z(n45626)) /* synthesis lut_function=(A (B (C+(D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam n728_bdd_3_lut_4_lut.init = 16'hf8f7;
    LUT4 i1_2_lut_rep_946_3_lut_4_lut (.A(n46110), .B(n46095), .C(n15_adj_316), 
         .D(n37_adj_301), .Z(n46067)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_946_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_125 (.A(n46110), .B(n46095), .C(n46090), 
         .D(n46136), .Z(n22924)) /* synthesis lut_function=(!((B (C (D)+!C !(D))+!B !(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_125.init = 16'h28a0;
    LUT4 i2_4_lut_adj_126 (.A(n160_adj_362), .B(n12_adj_395), .C(n161), 
         .D(n46039), .Z(n169)) /* synthesis lut_function=(!(A+(B (C)+!B (C+(D))))) */ ;
    defparam i2_4_lut_adj_126.init = 16'h0405;
    LUT4 n41402_bdd_4_lut (.A(n41402), .B(n41358), .C(n45898), .D(n45875), 
         .Z(n45566)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A !(((D)+!C)+!B))) */ ;
    defparam n41402_bdd_4_lut.init = 16'h5715;
    LUT4 i4555_2_lut_rep_757_3_lut_4_lut (.A(n46044), .B(n45892), .C(n4382[2]), 
         .D(n4382[1]), .Z(n45878)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i4555_2_lut_rep_757_3_lut_4_lut.init = 16'h0f2d;
    LUT4 mux_29_i5_3_lut (.A(n46852), .B(n46143), .C(n7), .Z(n112[4])) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_29_i5_3_lut.init = 16'hc5c5;
    LUT4 i2_4_lut_then_3_lut (.A(n23051), .B(n2046[5]), .C(n790[4]), .Z(n46867)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+!(C)))) */ ;
    defparam i2_4_lut_then_3_lut.init = 16'h6565;
    LUT4 i38121_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n46196), .B(n46048), 
         .C(n475[8]), .D(n45904), .Z(n43902)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (C))) */ ;
    defparam i38121_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0507;
    LUT4 i4557_2_lut_rep_758_3_lut_4_lut (.A(n46044), .B(n45892), .C(n4382[2]), 
         .D(n4382[1]), .Z(n45879)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i4557_2_lut_rep_758_3_lut_4_lut.init = 16'hf0d0;
    LUT4 i31574_1_lut_2_lut_3_lut_4_lut (.A(n46044), .B(n45892), .C(n4382[2]), 
         .D(n4382[1]), .Z(n38301)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A (C)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i31574_1_lut_2_lut_3_lut_4_lut.init = 16'hf0d2;
    LUT4 n338_bdd_4_lut (.A(n45845), .B(n330[2]), .C(n541[4]), .D(n45862), 
         .Z(n45571)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (C)) */ ;
    defparam n338_bdd_4_lut.init = 16'hf8d0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_127 (.A(n46110), .B(n46095), .C(n46136), 
         .D(n37_adj_301), .Z(n396[7])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_127.init = 16'h0080;
    LUT4 i1_3_lut_4_lut_adj_128 (.A(n45896), .B(n46124), .C(n45828), .D(n23030), 
         .Z(n4_adj_396)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;
    defparam i1_3_lut_4_lut_adj_128.init = 16'h7f80;
    LUT4 i15420_3_lut_rep_708_4_lut (.A(n45896), .B(n46124), .C(n1403[1]), 
         .D(n46145), .Z(n45829)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i15420_3_lut_rep_708_4_lut.init = 16'hf080;
    LUT4 i7251_2_lut_rep_944_3_lut_4_lut (.A(n124), .B(n46099), .C(n46088), 
         .D(n46143), .Z(n46065)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (B (C+(D))+!B (C))) */ ;
    defparam i7251_2_lut_rep_944_3_lut_4_lut.init = 16'hf6f0;
    CCU2D add_557_7 (.A0(n2345[4]), .B0(n2345[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40500), 
          .S0(n2358[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_557_7.INIT0 = 16'h5999;
    defparam add_557_7.INIT1 = 16'h0000;
    defparam add_557_7.INJECT1_0 = "NO";
    defparam add_557_7.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_129 (.A(n45756), .B(n45752), .C(n45740), .D(n30), 
         .Z(n2476[5])) /* synthesis lut_function=(!(A (B)+!A !(((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_4_lut_adj_129.init = 16'h7737;
    LUT4 div_28_i129_3_lut_4_lut (.A(n124), .B(n46099), .C(n46852), .D(n46143), 
         .Z(n23881)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D)))) */ ;
    defparam div_28_i129_3_lut_4_lut.init = 16'h9699;
    LUT4 mux_167_i4_4_lut (.A(n43701), .B(n46847), .C(n19), .D(n7_adj_397), 
         .Z(n755[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_167_i4_4_lut.init = 16'hcac5;
    LUT4 i2_4_lut_adj_130 (.A(n45636), .B(n45759), .C(n6_adj_398), .D(n45787), 
         .Z(n43701)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_4_lut_adj_130.init = 16'hd926;
    LUT4 i1_2_lut_rep_609_4_lut (.A(n23553), .B(n45733), .C(n44713), .Z(n45730)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_rep_609_4_lut.init = 16'h7878;
    LUT4 mux_1263_i1_4_lut (.A(n21510), .B(n4247[0]), .C(n46243), .D(n3611), 
         .Z(n3555[0])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(73[13] 82[22])
    defparam mux_1263_i1_4_lut.init = 16'hc0ca;
    LUT4 i2_2_lut_4_lut_3_lut_4_lut (.A(n45896), .B(n46124), .C(n45828), 
         .D(n1403[1]), .Z(n6_adj_399)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A ((D)+!C))) */ ;
    defparam i2_2_lut_4_lut_3_lut_4_lut.init = 16'h00f8;
    LUT4 i1_3_lut_rep_912_4_lut (.A(n16[8]), .B(n46100), .C(n43581), .D(n46041), 
         .Z(n46033)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_3_lut_rep_912_4_lut.init = 16'h8000;
    LUT4 mux_58_i6_3_lut_rep_866_4_lut (.A(n16[8]), .B(n46100), .C(n46179), 
         .D(n218[5]), .Z(n45987)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_58_i6_3_lut_rep_866_4_lut.init = 16'hf808;
    LUT4 i2_3_lut_4_lut_adj_131 (.A(n16[8]), .B(n46100), .C(n23650), .D(n43592), 
         .Z(n3[8])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i2_3_lut_4_lut_adj_131.init = 16'h0080;
    LUT4 n23541_bdd_4_lut (.A(n23541), .B(n45939), .C(n45919), .D(n45913), 
         .Z(n45585)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B (C+(D))+!B !(C+(D))))) */ ;
    defparam n23541_bdd_4_lut.init = 16'h399c;
    LUT4 i3_4_lut_adj_132 (.A(n22855), .B(n45968), .C(n8_adj_400), .D(n23445), 
         .Z(n43683)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i3_4_lut_adj_132.init = 16'h6996;
    LUT4 i2_3_lut_4_lut_adj_133 (.A(n45769), .B(n45786), .C(n45787), .D(n45761), 
         .Z(n7_adj_397)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_4_lut_adj_133.init = 16'hf708;
    LUT4 i2_3_lut_rep_679_4_lut (.A(n46051), .B(n45896), .C(n8_adj_401), 
         .D(n6_adj_402), .Z(n45800)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i2_3_lut_rep_679_4_lut.init = 16'hb44b;
    LUT4 i3993_2_lut_3_lut_4_lut (.A(n16[8]), .B(n46100), .C(n4_adj_403), 
         .D(n46055), .Z(n4233[3])) /* synthesis lut_function=(!(A (B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i3993_2_lut_3_lut_4_lut.init = 16'h7fff;
    LUT4 i1_2_lut_rep_762_3_lut_4_lut (.A(n46051), .B(n45896), .C(n545[8]), 
         .D(n46128), .Z(n45883)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_rep_762_3_lut_4_lut.init = 16'h78f0;
    LUT4 i15753_2_lut_3_lut_4_lut (.A(n16[8]), .B(n46100), .C(n4_adj_403), 
         .D(n46055), .Z(n22463)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i15753_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_125_i5_3_lut_4_lut (.A(n46051), .B(n45896), .C(n46128), .D(n1156[1]), 
         .Z(n545[4])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_125_i5_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_2_lut_rep_922_3_lut_4_lut (.A(n16[8]), .B(n46100), .C(n46055), 
         .D(n89_adj_303), .Z(n46043)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_922_3_lut_4_lut.init = 16'h0080;
    LUT4 i2046_2_lut_rep_760_3_lut_4_lut (.A(n46051), .B(n45896), .C(n545[8]), 
         .D(n46128), .Z(n45881)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2046_2_lut_rep_760_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i3818_3_lut_4_lut (.A(n46051), .B(n45896), .C(n45806), .D(n1156[1]), 
         .Z(n1169[2])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3818_3_lut_4_lut.init = 16'hf708;
    LUT4 i15131_2_lut_3_lut_4_lut (.A(n46051), .B(n45896), .C(n46137), 
         .D(n46115), .Z(n21753)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i15131_2_lut_3_lut_4_lut.init = 16'h6000;
    LUT4 i2_4_lut_adj_134 (.A(n46873), .B(oprand[2]), .C(n46878), .D(oprand[3]), 
         .Z(n30175)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;
    defparam i2_4_lut_adj_134.init = 16'h0444;
    LUT4 i1_3_lut (.A(oprand[3]), .B(oprand[2]), .C(oprand[4]), .Z(n87_adj_315)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i1_3_lut.init = 16'h2a2a;
    LUT4 i15027_4_lut (.A(n46090), .B(n15_adj_316), .C(n396[7]), .D(n46103), 
         .Z(n4330[1])) /* synthesis lut_function=(!(A ((C (D)+!C !(D))+!B)+!A !(B (C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i15027_4_lut.init = 16'h48c0;
    LUT4 i3_4_lut_4_lut_adj_135 (.A(n45725), .B(n45722), .C(n6_adj_404), 
         .D(n23094), .Z(n43707)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i3_4_lut_4_lut_adj_135.init = 16'h4bb4;
    LUT4 i2463_2_lut_3_lut_4_lut_4_lut (.A(n45899), .B(n45908), .C(n21[2]), 
         .D(n46848), .Z(n6574)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B+!(C (D))))) */ ;
    defparam i2463_2_lut_3_lut_4_lut_4_lut.init = 16'h1080;
    LUT4 i14937_3_lut_rep_752_4_lut_4_lut (.A(n45899), .B(n45908), .C(n21[2]), 
         .D(n46848), .Z(n45873)) /* synthesis lut_function=(A (B (C+(D)))+!A !(B+!(C+!(D)))) */ ;
    defparam i14937_3_lut_rep_752_4_lut_4_lut.init = 16'h9891;
    LUT4 n195_bdd_4_lut (.A(n45985), .B(n220_adj_405), .C(n45966), .D(n45941), 
         .Z(n45346)) /* synthesis lut_function=(A (B (C+(D))+!B (C+!(D)))+!A (B+!(C))) */ ;
    defparam n195_bdd_4_lut.init = 16'hede7;
    LUT4 i5_4_lut_rep_604 (.A(n44699), .B(n7_adj_406), .C(n45768), .D(n23553), 
         .Z(n45725)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i5_4_lut_rep_604.init = 16'h6996;
    LUT4 i2_2_lut_4_lut (.A(n45910), .B(n45899), .C(n45908), .D(n43759), 
         .Z(n6_adj_407)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (D))+!A !(B (C (D)+!C !(D))+!B (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_2_lut_4_lut.init = 16'h59a6;
    LUT4 i2437_4_lut_4_lut (.A(n45910), .B(n45908), .C(n45899), .D(n22852), 
         .Z(n6_adj_408)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A (B+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2437_4_lut_4_lut.init = 16'h20bb;
    LUT4 i1_2_lut_rep_954_3_lut_4_lut (.A(n46102), .B(n46118), .C(n37_adj_301), 
         .D(n46110), .Z(n46075)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_rep_954_3_lut_4_lut.init = 16'h0200;
    LUT4 i24038_2_lut_rep_956_3_lut_4_lut (.A(n46102), .B(n46118), .C(n46136), 
         .D(n46110), .Z(n46077)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i24038_2_lut_rep_956_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_3_lut_4_lut_adj_136 (.A(n45936), .B(n45901), .C(n43729), .D(n43768), 
         .Z(n41242)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i2_3_lut_4_lut_adj_136.init = 16'h6996;
    LUT4 i2_3_lut_4_lut_adj_137 (.A(n45900), .B(n45_adj_356), .C(n1156[2]), 
         .D(n46128), .Z(n4_adj_389)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i2_3_lut_4_lut_adj_137.init = 16'hfdff;
    LUT4 i2_2_lut_rep_960_3_lut_4_lut (.A(n46102), .B(n46118), .C(n23650), 
         .D(n46136), .Z(n46081)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i2_2_lut_rep_960_3_lut_4_lut.init = 16'h2000;
    LUT4 mux_132_i5_3_lut (.A(n1285[5]), .B(n545[4]), .C(n89_adj_320), 
         .Z(n1416[1])) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_132_i5_3_lut.init = 16'h5c5c;
    LUT4 i3056_3_lut_4_lut (.A(n45868), .B(n43686), .C(n45855), .D(n43675), 
         .Z(n8_adj_409)) /* synthesis lut_function=(A ((C (D))+!B)+!A !(B+!(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3056_3_lut_4_lut.init = 16'hb332;
    LUT4 n334_bdd_4_lut (.A(n45924), .B(n45877), .C(n46003), .D(n45865), 
         .Z(n45620)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C)+!B (C (D)+!C !(D))))) */ ;
    defparam n334_bdd_4_lut.init = 16'h2fbe;
    LUT4 i4115_2_lut_rep_706_3_lut_4_lut (.A(n45900), .B(n45_adj_356), .C(n1403[1]), 
         .D(n46124), .Z(n45827)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i4115_2_lut_rep_706_3_lut_4_lut.init = 16'h2000;
    LUT4 i14965_4_lut (.A(akku_o_c_0), .B(n4257[0]), .C(states_c[2]), 
         .D(data[0]), .Z(n21510)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(73[13] 82[22])
    defparam i14965_4_lut.init = 16'hc0c5;
    LUT4 mux_118_i5_3_lut (.A(n1012[5]), .B(n475[4]), .C(n45_adj_356), 
         .Z(n1156[1])) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_118_i5_3_lut.init = 16'h5c5c;
    CCU2D add_557_5 (.A0(n2345[2]), .B0(n2345[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2345[3]), .B1(n2345[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40499), .COUT(n40500), .S0(n2358[3]), .S1(n2358[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_557_5.INIT0 = 16'h5666;
    defparam add_557_5.INIT1 = 16'h5666;
    defparam add_557_5.INJECT1_0 = "NO";
    defparam add_557_5.INJECT1_1 = "NO";
    LUT4 mux_111_i5_4_lut (.A(n46086), .B(n462[4]), .C(n46196), .D(n46090), 
         .Z(n475[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_111_i5_4_lut.init = 16'hcac0;
    LUT4 i2_3_lut_rep_683_4_lut (.A(n45900), .B(n45_adj_356), .C(n46051), 
         .D(n6_adj_402), .Z(n45804)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C (D)))+!A (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i2_3_lut_rep_683_4_lut.init = 16'h0ff2;
    LUT4 i15377_2_lut_rep_950_3_lut_4_lut (.A(n16[8]), .B(n46106), .C(n46097), 
         .D(n46123), .Z(n46071)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i15377_2_lut_rep_950_3_lut_4_lut.init = 16'h8000;
    LUT4 i2_2_lut_3_lut_4_lut (.A(n45900), .B(n45_adj_356), .C(n46051), 
         .D(n6_adj_402), .Z(n6_adj_410)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i2_2_lut_3_lut_4_lut.init = 16'hf0f2;
    LUT4 i37177_3_lut_4_lut (.A(n16[8]), .B(n46106), .C(n46097), .D(n46109), 
         .Z(n23063)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)))+!A !(C (D)))) */ ;
    defparam i37177_3_lut_4_lut.init = 16'h7800;
    LUT4 i15095_3_lut_4_lut (.A(n45900), .B(n45_adj_356), .C(n1156[2]), 
         .D(n46128), .Z(n21696)) /* synthesis lut_function=(A (B (C (D))+!B !(C+!(D)))+!A (C (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i15095_3_lut_4_lut.init = 16'hd200;
    CCU2D add_557_3 (.A0(n2345[0]), .B0(n2345[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2345[1]), .B1(n2345[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40498), .COUT(n40499), .S0(n2358[1]), .S1(n2358[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_557_3.INIT0 = 16'h5666;
    defparam add_557_3.INIT1 = 16'h5999;
    defparam add_557_3.INJECT1_0 = "NO";
    defparam add_557_3.INJECT1_1 = "NO";
    CCU2D add_557_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n23806), .B1(n43670), .C1(n46138), .D1(n790[2]), .COUT(n40498), 
          .S1(n2358[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_557_1.INIT0 = 16'hF000;
    defparam add_557_1.INIT1 = 16'h06f6;
    defparam add_557_1.INJECT1_0 = "NO";
    defparam add_557_1.INJECT1_1 = "NO";
    CCU2D add_555_7 (.A0(n2332[4]), .B0(n2332[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40497), 
          .S0(n2345[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_555_7.INIT0 = 16'h5999;
    defparam add_555_7.INIT1 = 16'h0000;
    defparam add_555_7.INJECT1_0 = "NO";
    defparam add_555_7.INJECT1_1 = "NO";
    LUT4 mux_93_i6_3_lut_rep_742_4_lut (.A(n43686), .B(n45869), .C(n39_adj_343), 
         .D(n51_adj_344), .Z(n45863)) /* synthesis lut_function=(A (B+(C (D)))+!A !((C (D))+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_93_i6_3_lut_rep_742_4_lut.init = 16'haccc;
    LUT4 i4153_2_lut_rep_709_3_lut_4_lut (.A(n45900), .B(n45_adj_356), .C(n1403[1]), 
         .D(n46124), .Z(n45830)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i4153_2_lut_rep_709_3_lut_4_lut.init = 16'h2f0f;
    LUT4 i1_4_lut_rep_610_4_lut (.A(n45734), .B(n22479), .C(n2476[5]), 
         .D(n2476[2]), .Z(n45731)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A !(B (D)+!B !(C+!(D)))) */ ;
    defparam i1_4_lut_rep_610_4_lut.init = 16'h9a55;
    LUT4 n728_bdd_4_lut (.A(n720[1]), .B(n45763), .C(n45764), .D(n45770), 
         .Z(n45627)) /* synthesis lut_function=(A (B (C (D))+!B !(C+(D)))) */ ;
    defparam n728_bdd_4_lut.init = 16'h8002;
    LUT4 i1_2_lut_rep_940_3_lut_3_lut_4_lut_3_lut_4_lut (.A(n16[8]), .B(n46106), 
         .C(n46083), .D(n46097), .Z(n46061)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !((D)+!C))+!A !((D)+!C)) */ ;
    defparam i1_2_lut_rep_940_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h8078;
    LUT4 i2_4_lut_4_lut_adj_138 (.A(n2371[3]), .B(n2371[5]), .C(n6_adj_411), 
         .D(n2371[4]), .Z(n40779)) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_4_lut_4_lut_adj_138.init = 16'hdb24;
    LUT4 i15756_2_lut_3_lut_4_lut (.A(n45900), .B(n45_adj_356), .C(n1403[1]), 
         .D(n46124), .Z(n21707)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i15756_2_lut_3_lut_4_lut.init = 16'hf2f0;
    LUT4 mux_58_i4_3_lut (.A(n46064), .B(n218[3]), .C(n46179), .Z(n231_adj_515[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_58_i4_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_139 (.A(n45900), .B(n45_adj_356), .C(n8_adj_401), 
         .D(n46051), .Z(n5_adj_413)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_3_lut_4_lut_adj_139.init = 16'h0f2d;
    LUT4 div_46_i112_3_lut_rep_941_4_lut_3_lut_4_lut_3_lut_4_lut (.A(n16[8]), 
         .B(n46106), .C(n46083), .D(n46097), .Z(n46062)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+!(D)))+!A (C+!(D)))) */ ;
    defparam div_46_i112_3_lut_rep_941_4_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h0780;
    CCU2D add_555_5 (.A0(n2332[2]), .B0(n2332[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2332[3]), .B1(n2332[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40496), .COUT(n40497), .S0(n2345[3]), .S1(n2345[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_555_5.INIT0 = 16'h5666;
    defparam add_555_5.INIT1 = 16'h5666;
    defparam add_555_5.INJECT1_0 = "NO";
    defparam add_555_5.INJECT1_1 = "NO";
    FD1S3AX adreg_i2 (.D(adress_5__N_3[2]), .CK(clk_c), .Q(address[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam adreg_i2.GSR = "ENABLED";
    FD1S3AX adreg_i3 (.D(adress_5__N_3[3]), .CK(clk_c), .Q(address[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam adreg_i3.GSR = "ENABLED";
    FD1S3AX adreg_i4 (.D(adress_5__N_3[4]), .CK(clk_c), .Q(address[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam adreg_i4.GSR = "ENABLED";
    FD1S3AX adreg_i5 (.D(adress_5__N_3[5]), .CK(clk_c), .Q(address[5])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam adreg_i5.GSR = "ENABLED";
    FD1P3AX oprand_i0_i1 (.D(data[1]), .SP(clk_c_enable_26), .CK(clk_c), 
            .Q(oprand[1])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam oprand_i0_i1.GSR = "ENABLED";
    FD1P3AX oprand_i0_i2 (.D(data[2]), .SP(clk_c_enable_26), .CK(clk_c), 
            .Q(oprand[2])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam oprand_i0_i2.GSR = "ENABLED";
    FD1P3AX oprand_i0_i3 (.D(data[3]), .SP(clk_c_enable_26), .CK(clk_c), 
            .Q(oprand[3])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam oprand_i0_i3.GSR = "ENABLED";
    FD1P3AX oprand_i0_i4 (.D(data[4]), .SP(clk_c_enable_26), .CK(clk_c), 
            .Q(oprand[4])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam oprand_i0_i4.GSR = "ENABLED";
    FD1P3AX akku_i0_i2 (.D(n22540), .SP(clk_c_enable_22), .CK(clk_c), 
            .Q(akku_o_c_1)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam akku_i0_i2.GSR = "ENABLED";
    FD1P3AX akku_i0_i3 (.D(n22542), .SP(clk_c_enable_22), .CK(clk_c), 
            .Q(akku_o_c_2)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam akku_i0_i3.GSR = "ENABLED";
    FD1P3AX akku_i0_i4 (.D(n22544), .SP(clk_c_enable_22), .CK(clk_c), 
            .Q(akku_o_c_3)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam akku_i0_i4.GSR = "ENABLED";
    FD1P3AX akku_i0_i5 (.D(n22546), .SP(clk_c_enable_22), .CK(clk_c), 
            .Q(akku_o_c_4)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam akku_i0_i5.GSR = "ENABLED";
    FD1P3AX akku_i0_i6 (.D(n22548), .SP(clk_c_enable_22), .CK(clk_c), 
            .Q(akku_o_c_5)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam akku_i0_i6.GSR = "ENABLED";
    FD1P3AX akku_i0_i7 (.D(n3555[6]), .SP(clk_c_enable_22), .CK(clk_c), 
            .Q(akku_o_c_6)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam akku_i0_i7.GSR = "ENABLED";
    FD1P3AX akku_i0_i8 (.D(n3555[7]), .SP(clk_c_enable_22), .CK(clk_c), 
            .Q(akku_o_c_7)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam akku_i0_i8.GSR = "ENABLED";
    LUT4 i23888_2_lut_rep_765_3_lut_4_lut (.A(n45900), .B(n45_adj_356), 
         .C(n46128), .D(n46051), .Z(n45886)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i23888_2_lut_rep_765_3_lut_4_lut.init = 16'h2000;
    LUT4 i36947_2_lut_rep_764_3_lut_4_lut (.A(n45900), .B(n45_adj_356), 
         .C(n46115), .D(n46051), .Z(n45885)) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))+!A (C (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i36947_2_lut_rep_764_3_lut_4_lut.init = 16'hd020;
    LUT4 i14957_2_lut_3_lut_4_lut (.A(n45900), .B(n45_adj_356), .C(n46128), 
         .D(n46051), .Z(n4217[1])) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))+!A (C (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i14957_2_lut_3_lut_4_lut.init = 16'hd020;
    LUT4 i36917_2_lut_3_lut_4_lut (.A(n45900), .B(n45_adj_356), .C(n46122), 
         .D(n46051), .Z(n23019)) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))+!A (C (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i36917_2_lut_3_lut_4_lut.init = 16'hd020;
    LUT4 i2_4_lut_else_3_lut (.A(n23051), .B(n755[5]), .C(n755[6]), .D(n790[4]), 
         .Z(n46866)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !((C+!(D))+!B))) */ ;
    defparam i2_4_lut_else_3_lut.init = 16'h5955;
    LUT4 i15066_2_lut_rep_971_3_lut_4_lut (.A(n46136), .B(n46102), .C(n46106), 
         .D(n16[8]), .Z(n46092)) /* synthesis lut_function=(!(((C (D))+!B)+!A)) */ ;
    defparam i15066_2_lut_rep_971_3_lut_4_lut.init = 16'h0888;
    CCU2D add_555_3 (.A0(n2332[0]), .B0(n2332[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2332[1]), .B1(n2332[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40495), .COUT(n40496), .S0(n2345[1]), .S1(n2345[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_555_3.INIT0 = 16'h5666;
    defparam add_555_3.INIT1 = 16'h5999;
    defparam add_555_3.INJECT1_0 = "NO";
    defparam add_555_3.INJECT1_1 = "NO";
    CCU2D add_555_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n46870), .B1(n45750), .C1(n46146), .D1(n45757), .COUT(n40495), 
          .S1(n2345[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_555_1.INIT0 = 16'hF000;
    defparam add_555_1.INIT1 = 16'h04fe;
    defparam add_555_1.INJECT1_0 = "NO";
    defparam add_555_1.INJECT1_1 = "NO";
    CCU2D add_553_7 (.A0(n2319[4]), .B0(n2319[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40494), 
          .S0(n2332[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_553_7.INIT0 = 16'h5999;
    defparam add_553_7.INIT1 = 16'h0000;
    defparam add_553_7.INJECT1_0 = "NO";
    defparam add_553_7.INJECT1_1 = "NO";
    LUT4 i36941_2_lut_rep_972_3_lut_4_lut (.A(n46136), .B(n46102), .C(n46106), 
         .D(n16[8]), .Z(n46093)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(C (D)))) */ ;
    defparam i36941_2_lut_rep_972_3_lut_4_lut.init = 16'h7000;
    CCU2D add_553_5 (.A0(n2319[2]), .B0(n2319[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2319[3]), .B1(n2319[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40493), .COUT(n40494), .S0(n2332[3]), .S1(n2332[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_553_5.INIT0 = 16'h5666;
    defparam add_553_5.INIT1 = 16'h5666;
    defparam add_553_5.INJECT1_0 = "NO";
    defparam add_553_5.INJECT1_1 = "NO";
    CCU2D add_553_3 (.A0(n2319[0]), .B0(n2319[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2319[1]), .B1(n2319[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40492), .COUT(n40493), .S0(n2332[1]), .S1(n2332[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_553_3.INIT0 = 16'h5666;
    defparam add_553_3.INIT1 = 16'h5999;
    defparam add_553_3.INJECT1_0 = "NO";
    defparam add_553_3.INJECT1_1 = "NO";
    CCU2D add_553_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n46870), .B1(n2203[5]), .C1(n46146), .D1(n790[4]), .COUT(n40492), 
          .S1(n2332[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_553_1.INIT0 = 16'hF000;
    defparam add_553_1.INIT1 = 16'h04fe;
    defparam add_553_1.INJECT1_0 = "NO";
    defparam add_553_1.INJECT1_1 = "NO";
    FD1P3AX akku_i0_i9 (.D(n3555[8]), .SP(clk_c_enable_20), .CK(clk_c), 
            .Q(akku_o_c_8)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam akku_i0_i9.GSR = "ENABLED";
    LUT4 i24056_2_lut_3_lut_4_lut (.A(n15_adj_316), .B(n46103), .C(n46100), 
         .D(n37), .Z(n30783)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i24056_2_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_4_lut_adj_140 (.A(n45909), .B(n45903), .C(n231_adj_515[3]), 
         .D(n41358), .Z(n4_adj_384)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_140.init = 16'h9669;
    LUT4 div_39_i132_4_lut (.A(n160_adj_362), .B(n161), .C(n169), .D(n46023), 
         .Z(n190)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_i132_4_lut.init = 16'haaa9;
    LUT4 i15407_2_lut_rep_953_3_lut_4_lut (.A(n15_adj_316), .B(n46103), 
         .C(n46196), .D(n37), .Z(n46074)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i15407_2_lut_rep_953_3_lut_4_lut.init = 16'h0080;
    LUT4 i7241_2_lut_rep_952_3_lut_4_lut (.A(n46112), .B(n46143), .C(n124), 
         .Z(n46073)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i7241_2_lut_rep_952_3_lut_4_lut.init = 16'h4848;
    LUT4 mux_29_i6_3_lut_4_lut (.A(n46112), .B(n7), .C(n124), .Z(n112[5])) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_29_i6_3_lut_4_lut.init = 16'he2e2;
    LUT4 i2_3_lut_4_lut_adj_141 (.A(n45903), .B(n45909), .C(n231_adj_515[3]), 
         .D(n40830), .Z(n41402)) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_4_lut_adj_141.init = 16'hdb24;
    LUT4 i1961_4_lut_3_lut_4_lut (.A(n45903), .B(n45909), .C(n231_adj_515[3]), 
         .D(n40830), .Z(n6_adj_414)) /* synthesis lut_function=(A (B+!(C (D)))+!A !((C+(D))+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1961_4_lut_3_lut_4_lut.init = 16'h8aae;
    LUT4 i1_2_lut_rep_773_4_lut (.A(n45903), .B(n231_adj_515[3]), .C(n37_adj_318), 
         .D(n45908), .Z(n45894)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_773_4_lut.init = 16'h53ac;
    LUT4 i23840_2_lut_3_lut_4_lut (.A(n46112), .B(n46143), .C(n124), .Z(n12_adj_358)) /* synthesis lut_function=(A ((C)+!B)+!A !(B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i23840_2_lut_3_lut_4_lut.init = 16'hb7b7;
    LUT4 i1_2_lut_rep_955_3_lut_4_lut (.A(n46118), .B(n46106), .C(n46110), 
         .D(n16[8]), .Z(n46076)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_2_lut_rep_955_3_lut_4_lut.init = 16'h4000;
    LUT4 n22905_bdd_4_lut (.A(n6_adj_398), .B(n45764), .C(n45759), .D(n1947[2]), 
         .Z(n45632)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B ((D)+!C)+!B !(C (D))))) */ ;
    defparam n22905_bdd_4_lut.init = 16'h32c8;
    LUT4 i24233_2_lut_rep_766_3_lut_4_lut (.A(n45904), .B(n46196), .C(n46122), 
         .D(n45_adj_356), .Z(n45887)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i24233_2_lut_rep_766_3_lut_4_lut.init = 16'h0080;
    LUT4 i24236_2_lut_rep_767_3_lut_4_lut (.A(n45904), .B(n46196), .C(n46124), 
         .D(n45_adj_356), .Z(n45888)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i24236_2_lut_rep_767_3_lut_4_lut.init = 16'h0080;
    LUT4 mux_40_i7_3_lut_rep_962_4_lut_4_lut (.A(n46107), .B(n102), .C(n11), 
         .D(n67), .Z(n46083)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_40_i7_3_lut_rep_962_4_lut_4_lut.init = 16'hcec0;
    LUT4 i6781_2_lut_rep_948_4_lut_4_lut_4_lut (.A(n46107), .B(n102), .C(n67), 
         .D(n46078), .Z(n46069)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i6781_2_lut_rep_948_4_lut_4_lut_4_lut.init = 16'h8a08;
    LUT4 i15139_2_lut_rep_643_3_lut_4_lut (.A(n46847), .B(n45788), .C(n45787), 
         .D(n45786), .Z(n45764)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i15139_2_lut_rep_643_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_2_lut_rep_966_3_lut_4_lut (.A(n46108), .B(n46121), .C(n46110), 
         .D(n46118), .Z(n46087)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_2_lut_rep_966_3_lut_4_lut.init = 16'h0080;
    LUT4 i23778_2_lut_rep_768_3_lut_4_lut (.A(n45904), .B(n46196), .C(n46115), 
         .D(n45_adj_356), .Z(n45889)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i23778_2_lut_rep_768_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_963_3_lut_4_lut (.A(n46108), .B(n46121), .C(n46123), 
         .D(n46136), .Z(n46084)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_963_3_lut_4_lut.init = 16'h8000;
    LUT4 n6_bdd_4_lut (.A(n45764), .B(n45763), .C(n45759), .D(n1947[2]), 
         .Z(n45634)) /* synthesis lut_function=(A (C (D))+!A !(B ((D)+!C)+!B !(C (D)))) */ ;
    defparam n6_bdd_4_lut.init = 16'hb040;
    LUT4 i15067_2_lut_rep_769_3_lut_4_lut (.A(n45904), .B(n46196), .C(n46051), 
         .D(n45_adj_356), .Z(n45890)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i15067_2_lut_rep_769_3_lut_4_lut.init = 16'hfff7;
    LUT4 i3799_2_lut_rep_770_3_lut_4_lut (.A(n45904), .B(n46196), .C(n46051), 
         .D(n45_adj_356), .Z(n45891)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i3799_2_lut_rep_770_3_lut_4_lut.init = 16'h0080;
    LUT4 i23777_2_lut_rep_771_3_lut_4_lut (.A(n45904), .B(n46196), .C(n46111), 
         .D(n45_adj_356), .Z(n45892)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i23777_2_lut_rep_771_3_lut_4_lut.init = 16'h0080;
    LUT4 i4537_1_lut_2_lut_3_lut_4_lut (.A(n45904), .B(n46196), .C(n46111), 
         .D(n45_adj_356), .Z(n4400[0])) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i4537_1_lut_2_lut_3_lut_4_lut.init = 16'hff7f;
    LUT4 i24117_2_lut_rep_961_3_lut_4_lut (.A(n46108), .B(n46121), .C(n46136), 
         .D(n46118), .Z(n46082)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i24117_2_lut_rep_961_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_964_3_lut_4_lut (.A(n46108), .B(n46121), .C(n46109), 
         .D(n46136), .Z(n46085)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_964_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_142 (.A(n45919), .B(n41244), .C(n45913), .D(n23541), 
         .Z(n5_adj_415)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A !(B+!((D)+!C)))) */ ;
    defparam i1_4_lut_adj_142.init = 16'h6e76;
    LUT4 i15405_2_lut_rep_965_3_lut_4_lut (.A(n37_adj_301), .B(n46110), 
         .C(n37), .D(n15_adj_316), .Z(n46086)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i15405_2_lut_rep_965_3_lut_4_lut.init = 16'h0400;
    LUT4 i2_3_lut_adj_143 (.A(n45947), .B(n22855), .C(n45987), .Z(n23541)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i2_3_lut_adj_143.init = 16'h9696;
    LUT4 i2_4_lut_adj_144 (.A(n43785), .B(n405[2]), .C(n6734), .D(n6_adj_416), 
         .Z(n43729)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B (D)+!B !(D))) */ ;
    defparam i2_4_lut_adj_144.init = 16'hc639;
    LUT4 i36915_4_lut (.A(n22902), .B(n45880), .C(n22900), .D(n45876), 
         .Z(n43785)) /* synthesis lut_function=(A+!(((D)+!C)+!B)) */ ;
    defparam i36915_4_lut.init = 16'haaea;
    LUT4 i2_3_lut_adj_145 (.A(n3[4]), .B(n45929), .C(n45940), .Z(n22900)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i2_3_lut_adj_145.init = 16'h9696;
    LUT4 n1147_bdd_4_lut_38385 (.A(n45896), .B(n46051), .C(n46128), .D(n1156[2]), 
         .Z(n45652)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C)))) */ ;
    defparam n1147_bdd_4_lut_38385.init = 16'h6040;
    LUT4 mux_58_i2_3_lut_rep_781 (.A(n218[4]), .B(n218[1]), .C(n46179), 
         .Z(n45902)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_58_i2_3_lut_rep_781.init = 16'hcaca;
    LUT4 mux_40_i6_3_lut_rep_921_4_lut (.A(n46069), .B(n130_adj_360), .C(n11), 
         .D(n46078), .Z(n46042)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_40_i6_3_lut_rep_921_4_lut.init = 16'hfe0e;
    LUT4 n45635_bdd_3_lut_4_lut (.A(n46847), .B(n45788), .C(n45632), .D(n45635), 
         .Z(n45636)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam n45635_bdd_3_lut_4_lut.init = 16'hf960;
    LUT4 i2_4_lut_adj_146 (.A(n8_adj_409), .B(n22924), .C(n45918), .D(n4_adj_417), 
         .Z(n40941)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i2_4_lut_adj_146.init = 16'h6996;
    LUT4 mux_65_i4_3_lut_rep_778_4_lut (.A(n22855), .B(n45905), .C(n37_adj_318), 
         .D(n231_adj_515[3]), .Z(n45899)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_65_i4_3_lut_rep_778_4_lut.init = 16'h6f60;
    LUT4 akku_o_c_0_bdd_4_lut (.A(akku_o_c_0), .B(akku_o_c_3), .C(akku_o_c_4), 
         .D(akku_o_c_1), .Z(n46869)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;
    defparam akku_o_c_0_bdd_4_lut.init = 16'h9009;
    LUT4 i3_4_lut_adj_147 (.A(n45906), .B(n4_adj_418), .C(n6_adj_419), 
         .D(n8_adj_420), .Z(n43714)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i3_4_lut_adj_147.init = 16'h6996;
    LUT4 i1_4_lut_4_lut_adj_148 (.A(n22855), .B(n45905), .C(n6_adj_414), 
         .D(n22867), .Z(n7_adj_421)) /* synthesis lut_function=(!(A (B (C+!(D))+!B ((D)+!C))+!A !(B ((D)+!C)+!B (C+!(D))))) */ ;
    defparam i1_4_lut_4_lut_adj_148.init = 16'h5c35;
    LUT4 i2_3_lut_rep_777_4_lut (.A(n22855), .B(n45905), .C(n231_adj_515[3]), 
         .D(n45909), .Z(n45898)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i2_3_lut_rep_777_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_969_3_lut_4_lut (.A(n46120), .B(n46108), .C(n16[8]), 
         .D(n46118), .Z(n46090)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_969_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_adj_149 (.A(n43695), .B(n43750), .Z(n41286)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_149.init = 16'h6666;
    LUT4 i1_2_lut_2_lut (.A(n45774), .B(n6_adj_422), .Z(n40913)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut_2_lut.init = 16'h9999;
    LUT4 i3_4_lut_adj_150 (.A(n8_adj_423), .B(n45854), .C(n40941), .D(n43675), 
         .Z(n41291)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i3_4_lut_adj_150.init = 16'h6996;
    LUT4 i2_2_lut_3_lut (.A(n22855), .B(n45905), .C(n41358), .Z(n7_adj_424)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i2_2_lut_3_lut.init = 16'h9696;
    LUT4 n271_bdd_4_lut_38352 (.A(n270_adj_516[6]), .B(n270_adj_516[5]), 
         .C(n270_adj_516[3]), .D(n270_adj_516[4]), .Z(n45348)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n271_bdd_4_lut_38352.init = 16'hfffe;
    LUT4 i1_2_lut_rep_968_3_lut_3_lut_4_lut (.A(n46207), .B(n46113), .C(n67), 
         .D(n102), .Z(n46089)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (C+!(D)))) */ ;
    defparam i1_2_lut_rep_968_3_lut_3_lut_4_lut.init = 16'h0f80;
    LUT4 n1147_bdd_4_lut (.A(n45896), .B(n46051), .C(n46128), .D(n1156[2]), 
         .Z(n45653)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C (D)))+!A !(B (C))) */ ;
    defparam n1147_bdd_4_lut.init = 16'h9f3f;
    LUT4 i1_2_lut_rep_980_4_lut (.A(n46207), .B(n46113), .C(n67), .D(n102), 
         .Z(n46101)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i1_2_lut_rep_980_4_lut.init = 16'hf080;
    LUT4 i24505_2_lut_3_lut_4_lut (.A(n46207), .B(n46113), .C(n67), .D(n102), 
         .Z(n130_adj_360)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;
    defparam i24505_2_lut_3_lut_4_lut.init = 16'h0070;
    LUT4 div_39_i91_3_lut_rep_970_4_lut_3_lut_4_lut (.A(n46207), .B(n46113), 
         .C(n67), .D(n102), .Z(n46091)) /* synthesis lut_function=(A (B ((D)+!C))) */ ;
    defparam div_39_i91_3_lut_rep_970_4_lut_3_lut_4_lut.init = 16'h8808;
    LUT4 n276_bdd_4_lut_38390 (.A(n270[3]), .B(n270[8]), .C(n270[4]), 
         .D(n270[7]), .Z(n45661)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n276_bdd_4_lut_38390.init = 16'hfffe;
    LUT4 i1_2_lut_rep_975_3_lut_4_lut (.A(n46207), .B(n11), .C(n16[8]), 
         .D(n46120), .Z(n46096)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_975_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_151 (.A(n46179), .B(n46064), .C(n23063), 
         .D(n46085), .Z(n23445)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_151.init = 16'hf078;
    LUT4 n276_bdd_4_lut (.A(n255), .B(n251), .C(n254), .D(n250), .Z(n45662)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n276_bdd_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_adj_152 (.A(n45856), .B(n43686), .C(n45869), .Z(n640[1])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;
    defparam i2_3_lut_adj_152.init = 16'h6969;
    LUT4 i1_2_lut_rep_976_3_lut_4_lut (.A(n46207), .B(n11), .C(n46136), 
         .D(n46121), .Z(n46097)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_976_3_lut_4_lut.init = 16'h8000;
    LUT4 i23864_2_lut_rep_779_4_lut (.A(n45906), .B(n45914), .C(n37), 
         .D(n46196), .Z(n45900)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (D)+!B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i23864_2_lut_rep_779_4_lut.init = 16'h5c00;
    LUT4 i1_2_lut_rep_974_3_lut_4_lut (.A(n46207), .B(n11), .C(n46118), 
         .D(n46121), .Z(n46095)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_974_3_lut_4_lut.init = 16'h0800;
    LUT4 i2_2_lut_rep_979_3_lut_4_lut (.A(n46207), .B(n11), .C(n46118), 
         .D(n46120), .Z(n46100)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i2_2_lut_rep_979_3_lut_4_lut.init = 16'h0800;
    LUT4 i2575_3_lut_rep_780_3_lut (.A(n45940), .B(n45929), .C(n3[4]), 
         .Z(n45901)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2575_3_lut_rep_780_3_lut.init = 16'hd4d4;
    LUT4 n45346_bdd_4_lut_38353 (.A(n251_adj_429), .B(n45956), .C(n254_adj_430), 
         .D(n45950), .Z(n45351)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n45346_bdd_4_lut_38353.init = 16'hfffe;
    LUT4 n45351_bdd_2_lut (.A(n45351), .B(n45346), .Z(n45352)) /* synthesis lut_function=(A+(B)) */ ;
    defparam n45351_bdd_2_lut.init = 16'heeee;
    LUT4 i4639_2_lut_rep_648_4_lut (.A(n1829[5]), .B(n685[3]), .C(n89), 
         .D(n45788), .Z(n45769)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B (D)+!B ((D)+!C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i4639_2_lut_rep_648_4_lut.init = 16'h005c;
    LUT4 i1_2_lut_rep_933_3_lut_4_lut_4_lut (.A(n46179), .B(n46118), .C(n46064), 
         .D(n46097), .Z(n46054)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))) */ ;
    defparam i1_2_lut_rep_933_3_lut_4_lut_4_lut.init = 16'h82a0;
    LUT4 i2234_2_lut_rep_925_3_lut_4_lut_4_lut (.A(n46179), .B(n46118), 
         .C(n46064), .D(n46097), .Z(n46046)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))) */ ;
    defparam i2234_2_lut_rep_925_3_lut_4_lut_4_lut.init = 16'h80a0;
    LUT4 i3_4_lut_adj_153 (.A(n21418), .B(n6_adj_431), .C(n4_adj_363), 
         .D(n45874), .Z(n583)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3_4_lut_adj_153.init = 16'h6996;
    LUT4 i2_4_lut_adj_154 (.A(n21482), .B(n43689), .C(n541[4]), .D(n45862), 
         .Z(n6_adj_431)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))+!B !(C+(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_4_lut_adj_154.init = 16'h6663;
    LUT4 i14946_4_lut (.A(n23447), .B(n541[4]), .C(n330[2]), .D(n45862), 
         .Z(n21482)) /* synthesis lut_function=(!(A+(B ((D)+!C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i14946_4_lut.init = 16'h1151;
    LUT4 i1_2_lut_rep_982_4_lut (.A(n46114), .B(n15), .C(n23650), .D(n37_adj_301), 
         .Z(n46103)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_982_4_lut.init = 16'h0040;
    LUT4 i3_3_lut_rep_784 (.A(n5_adj_415), .B(n23515), .C(n45928), .Z(n45905)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i3_3_lut_rep_784.init = 16'h9696;
    LUT4 i5584_4_lut_4_lut (.A(n2629[2]), .B(n2629[5]), .C(n2629[1]), 
         .D(n2_adj_367), .Z(n6_adj_432)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5584_4_lut_4_lut.init = 16'hecc8;
    LUT4 i1_2_lut_rep_782_4_lut (.A(n5_adj_415), .B(n23515), .C(n45928), 
         .D(n22855), .Z(n45903)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i1_2_lut_rep_782_4_lut.init = 16'h6996;
    LUT4 i37290_2_lut_rep_978_3_lut_4_lut (.A(n46116), .B(n124), .C(n46117), 
         .Z(n46099)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i37290_2_lut_rep_978_3_lut_4_lut.init = 16'hf8f8;
    LUT4 mux_107_i7_3_lut_rep_783_4_lut (.A(n22635), .B(n45907), .C(n37), 
         .D(n45914), .Z(n45904)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_107_i7_3_lut_rep_783_4_lut.init = 16'h1f10;
    LUT4 i1_4_lut_adj_155 (.A(n8_adj_433), .B(n45871), .C(n45880), .D(n45876), 
         .Z(n43768)) /* synthesis lut_function=(!(A (B+(C (D)))+!A !(B+(C (D))))) */ ;
    defparam i1_4_lut_adj_155.init = 16'h5666;
    LUT4 i2_3_lut_4_lut_adj_156 (.A(n22635), .B(n45907), .C(n45914), .D(n45859), 
         .Z(n22978)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_4_lut_adj_156.init = 16'he11e;
    LUT4 mux_58_i3_3_lut_rep_788 (.A(n218[5]), .B(n218[2]), .C(n46179), 
         .Z(n45909)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_58_i3_3_lut_rep_788.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_157 (.A(n218[5]), .B(n218[2]), .C(n46179), 
         .D(n41358), .Z(n4_adj_357)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_4_lut_adj_157.init = 16'h35ca;
    LUT4 mux_65_i3_3_lut (.A(n41358), .B(n45909), .C(n37_adj_318), .Z(n21[2])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_65_i3_3_lut.init = 16'hacac;
    LUT4 div_28_i106_3_lut_4_lut_3_lut_4_lut (.A(n46116), .B(n124), .C(n46117), 
         .Z(n152)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_i106_3_lut_4_lut_3_lut_4_lut.init = 16'h8080;
    LUT4 i5_4_lut (.A(n43683), .B(n7_adj_421), .C(n45976), .D(n45585), 
         .Z(n41358)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i5_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_649_4_lut (.A(n1829[5]), .B(n685[3]), .C(n89), .D(n45788), 
         .Z(n45770)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(B (D)+!B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_649_4_lut.init = 16'ha35c;
    LUT4 i23735_4_lut (.A(n40779), .B(n46157), .C(n825[0]), .D(n45), 
         .Z(n895[0])) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i23735_4_lut.init = 16'h88c0;
    PFUMX i38229 (.BLUT(n45352), .ALUT(n45350), .C0(n45930), .Z(n43333));
    LUT4 div_28_i107_3_lut_rep_967_4_lut_4_lut (.A(n46116), .B(n124), .C(n46117), 
         .Z(n46088)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_i107_3_lut_rep_967_4_lut_4_lut.init = 16'h6262;
    LUT4 i15204_3_lut_rep_611_4_lut (.A(n45747), .B(n45736), .C(n23553), 
         .Z(n45732)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i15204_3_lut_rep_611_4_lut.init = 16'he0e0;
    LUT4 i14939_3_lut_rep_774_4_lut (.A(n45915), .B(n46012), .C(n45899), 
         .D(n45908), .Z(n45895)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(B (C+(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i14939_3_lut_rep_774_4_lut.init = 16'h6660;
    LUT4 mux_33_i6_3_lut_rep_957_4_lut (.A(n46136), .B(n46121), .C(n46207), 
         .D(n112[5]), .Z(n46078)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam mux_33_i6_3_lut_rep_957_4_lut.init = 16'hf808;
    LUT4 i23817_2_lut_3_lut_4_lut (.A(n46069), .B(n130_adj_360), .C(n46050), 
         .D(n46078), .Z(n12_adj_395)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B (C+(D))))) */ ;
    defparam i23817_2_lut_3_lut_4_lut.init = 16'h0e01;
    LUT4 i2_3_lut_4_lut_4_lut_adj_158 (.A(n46059), .B(n45914), .C(n45859), 
         .D(n45906), .Z(n41108)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !((D)+!C))+!A !(B (C+!(D))+!B !((D)+!C)))) */ ;
    defparam i2_3_lut_4_lut_4_lut_adj_158.init = 16'h6a56;
    LUT4 i3470_4_lut_3_lut_4_lut_4_lut (.A(n46059), .B(n45914), .C(n45859), 
         .D(n45906), .Z(n6_adj_419)) /* synthesis lut_function=(A (B (C (D))+!B (C+(D)))+!A (D)) */ ;
    defparam i3470_4_lut_3_lut_4_lut_4_lut.init = 16'hf720;
    LUT4 i4_4_lut_adj_159 (.A(n213), .B(n211), .C(n215), .D(n6_adj_300), 
         .Z(n22716)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i4_4_lut_adj_159.init = 16'hfffe;
    LUT4 i2_3_lut_rep_989_4_lut (.A(n43592), .B(n37_adj_340), .C(n23650), 
         .D(n15), .Z(n46110)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_3_lut_rep_989_4_lut.init = 16'h1000;
    LUT4 i3441_2_lut_rep_785_3_lut_4_lut (.A(n46059), .B(n45914), .C(n22635), 
         .D(n4330[1]), .Z(n45906)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3441_2_lut_rep_785_3_lut_4_lut.init = 16'hfffd;
    LUT4 i1_2_lut_rep_700_3_lut_4_lut_4_lut (.A(n46122), .B(n89_adj_303), 
         .C(n45829), .D(n45896), .Z(n45821)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A (B+!(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_700_3_lut_4_lut_4_lut.init = 16'h1230;
    LUT4 i1_2_lut_rep_983_3_lut_4_lut (.A(n46122), .B(n89_adj_303), .C(n43547), 
         .D(n46137), .Z(n46104)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_983_3_lut_4_lut.init = 16'h2000;
    LUT4 i2_2_lut_4_lut_adj_160 (.A(n222_adj_334), .B(n20[6]), .C(n45916), 
         .D(n253), .Z(n8_adj_434)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_2_lut_4_lut_adj_160.init = 16'hffca;
    LUT4 i2_3_lut_4_lut_adj_161 (.A(n45919), .B(n231_adj_515[3]), .C(n45947), 
         .D(n23541), .Z(n22867)) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_4_lut_adj_161.init = 16'hdb24;
    LUT4 mux_111_i3_3_lut_4_lut (.A(n45917), .B(n15_adj_316), .C(n46196), 
         .D(n462[2]), .Z(n475[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_111_i3_3_lut_4_lut.init = 16'hf808;
    LUT4 i14916_3_lut_rep_739_4_lut_4_lut (.A(n3[3]), .B(n45866), .C(n3[2]), 
         .D(n427[1]), .Z(n45860)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i14916_3_lut_rep_739_4_lut_4_lut.init = 16'hf700;
    LUT4 i3_4_lut_adj_162 (.A(n45973), .B(n221_adj_435), .C(n45972), .D(n220_adj_405), 
         .Z(n22712)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3_4_lut_adj_162.init = 16'hffdf;
    LUT4 i1_2_lut_3_lut_4_lut_adj_163 (.A(n45917), .B(n15_adj_316), .C(n4330[1]), 
         .D(n46059), .Z(n4_adj_418)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_3_lut_4_lut_adj_163.init = 16'h780f;
    LUT4 i3434_2_lut_rep_786_3_lut_4_lut (.A(n45917), .B(n15_adj_316), .C(n4330[1]), 
         .D(n46059), .Z(n45907)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (C+!(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i3434_2_lut_rep_786_3_lut_4_lut.init = 16'hf8ff;
    LUT4 i3_4_lut_rep_653 (.A(n45775), .B(n6_adj_376), .C(n23779), .D(n45792), 
         .Z(n45774)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i3_4_lut_rep_653.init = 16'h6996;
    LUT4 i2389_2_lut_rep_789_4_lut (.A(n45919), .B(n45947), .C(n37_adj_318), 
         .D(n46012), .Z(n45910)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i2389_2_lut_rep_789_4_lut.init = 16'h53ac;
    LUT4 div_53_i176_3_lut_rep_791_4_lut (.A(n45922), .B(n22673), .C(n20[6]), 
         .D(n222_adj_334), .Z(n45912)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_i176_3_lut_rep_791_4_lut.init = 16'hf1e0;
    LUT4 div_53_i177_3_lut_4_lut (.A(n45922), .B(n22673), .C(n20[5]), 
         .D(n223), .Z(n253)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_i177_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i38391 (.BLUT(n45662), .ALUT(n45661), .C0(n208[1]), .Z(n45663));
    LUT4 div_53_i179_3_lut_4_lut (.A(n45922), .B(n22673), .C(n20[3]), 
         .D(n45926), .Z(n255)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_i179_3_lut_4_lut.init = 16'he0f1;
    LUT4 mux_54_i3_3_lut_4_lut (.A(n45922), .B(n22673), .C(n29_adj_353), 
         .D(n73_adj_336), .Z(n218[2])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_54_i3_3_lut_4_lut.init = 16'hefe0;
    LUT4 div_53_i174_3_lut_4_lut (.A(n45922), .B(n22673), .C(n20[8]), 
         .D(n220), .Z(n250)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_i174_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_53_i180_3_lut_4_lut (.A(n45922), .B(n22673), .C(n20[2]), 
         .D(n73_adj_336), .Z(n256)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_i180_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_53_i178_3_lut_4_lut (.A(n45922), .B(n22673), .C(n20[4]), 
         .D(n45925), .Z(n254)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_i178_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_53_i175_3_lut_4_lut (.A(n45922), .B(n22673), .C(n20[7]), 
         .D(n221_adj_333), .Z(n251)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_i175_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3427_2_lut_rep_790_3_lut_4_lut (.A(n45923), .B(n37_adj_301), .C(n46059), 
         .D(n15_adj_316), .Z(n45911)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i3427_2_lut_rep_790_3_lut_4_lut.init = 16'h2f0f;
    LUT4 i1_2_lut_4_lut_adj_164 (.A(n40740), .B(n45782), .C(n6_adj_422), 
         .D(n6_adj_376), .Z(n5_adj_436)) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_4_lut_adj_164.init = 16'h8e71;
    LUT4 i3_4_lut_adj_165 (.A(n223), .B(n220), .C(n221_adj_333), .D(n222_adj_334), 
         .Z(n22673)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3_4_lut_adj_165.init = 16'hfffe;
    LUT4 i3210_2_lut_4_lut_4_lut (.A(n45923), .B(n37_adj_301), .C(n45869), 
         .D(n43686), .Z(n754[2])) /* synthesis lut_function=(A (B (D)+!B !(C))+!A (B (D)+!B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i3210_2_lut_4_lut_4_lut.init = 16'hde12;
    LUT4 i2_3_lut_4_lut_adj_166 (.A(n46870), .B(n7), .C(n46207), .D(n16[8]), 
         .Z(n67)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_3_lut_4_lut_adj_166.init = 16'h8000;
    LUT4 i2_3_lut_4_lut_4_lut_adj_167 (.A(n46085), .B(n46056), .C(n45987), 
         .D(n46027), .Z(n23515)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C+(D))+!B (C (D)))) */ ;
    defparam i2_3_lut_4_lut_4_lut_adj_167.init = 16'ha995;
    LUT4 i1_2_lut_rep_985_3_lut_4_lut (.A(n46870), .B(n7), .C(n11), .D(n46207), 
         .Z(n46106)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_985_3_lut_4_lut.init = 16'h8000;
    LUT4 i63_then_4_lut_adj_168 (.A(akku_o_c_0), .B(n46189), .C(n117_adj_323), 
         .D(n122_adj_437), .Z(n46294)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i63_then_4_lut_adj_168.init = 16'h8000;
    LUT4 n398_bdd_3_lut_rep_740_4_lut (.A(n45923), .B(n37_adj_301), .C(n45863), 
         .D(n396[7]), .Z(n45861)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam n398_bdd_3_lut_rep_740_4_lut.init = 16'hdfff;
    LUT4 n6_bdd_4_lut_4_lut (.A(n46077), .B(n45923), .C(n45869), .D(n46076), 
         .Z(n43686)) /* synthesis lut_function=(A (B (D)+!B (C (D)))) */ ;
    defparam n6_bdd_4_lut_4_lut.init = 16'ha800;
    LUT4 i2_3_lut_4_lut_adj_169 (.A(n46027), .B(n43683), .C(n45947), .D(n231_adj_515[3]), 
         .Z(n40830)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i2_3_lut_4_lut_adj_169.init = 16'h6996;
    LUT4 i2_4_lut_adj_170 (.A(n45583), .B(n45895), .C(n6574), .D(n22852), 
         .Z(n43759)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_4_lut_adj_170.init = 16'hc936;
    LUT4 i1_4_lut_adj_171 (.A(n15_adj_438), .B(n3622), .C(n13), .D(n14_adj_439), 
         .Z(n4_adj_440)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_171.init = 16'hccc8;
    LUT4 i2129_4_lut_3_lut_rep_792_4_lut (.A(n46027), .B(n43683), .C(n45947), 
         .D(n231_adj_515[3]), .Z(n45913)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C+!(D))))) */ ;
    defparam i2129_4_lut_3_lut_rep_792_4_lut.init = 16'h6f06;
    LUT4 i2_2_lut_rep_986_3_lut_4_lut (.A(n46132), .B(n7), .C(n46207), 
         .D(n46136), .Z(n46107)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i2_2_lut_rep_986_3_lut_4_lut.init = 16'he000;
    LUT4 i1_2_lut_rep_981_3_lut_4_lut (.A(n46132), .B(n7), .C(n11), .D(n46207), 
         .Z(n46102)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_981_3_lut_4_lut.init = 16'he000;
    LUT4 i17149_2_lut_rep_990_3_lut_4_lut (.A(n46145), .B(n46124), .C(n46137), 
         .D(n89_adj_303), .Z(n46111)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i17149_2_lut_rep_990_3_lut_4_lut.init = 16'h0080;
    LUT4 i621_1_lut_3_lut_4_lut (.A(n46130), .B(n45778), .C(n23081), .D(n43991), 
         .Z(n2662)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B+((D)+!C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i621_1_lut_3_lut_4_lut.init = 16'h00b0;
    LUT4 i2_3_lut_rep_652_4_lut (.A(n46130), .B(n45778), .C(n23081), .D(n43991), 
         .Z(n45773)) /* synthesis lut_function=(A ((D)+!C)+!A (B+((D)+!C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_rep_652_4_lut.init = 16'hff4f;
    LUT4 mux_65_i5_3_lut_rep_794_4_lut (.A(n46027), .B(n43683), .C(n37_adj_318), 
         .D(n45947), .Z(n45915)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_65_i5_3_lut_rep_794_4_lut.init = 16'h6f60;
    LUT4 i2_4_lut_adj_172 (.A(n41108), .B(n45834), .C(n21624), .D(n7658), 
         .Z(n43762)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+(D)))) */ ;
    defparam i2_4_lut_adj_172.init = 16'h9996;
    LUT4 n45395_bdd_4_lut (.A(n46261), .B(n46266), .C(n46882), .D(akku_o_c_2), 
         .Z(n45691)) /* synthesis lut_function=(!(A+(B (C+(D))+!B (C+!(D))))) */ ;
    defparam n45395_bdd_4_lut.init = 16'h0104;
    LUT4 mux_29_i7_3_lut_4_lut_4_lut (.A(n46125), .B(n93), .C(n7), .D(n46126), 
         .Z(n112[6])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_29_i7_3_lut_4_lut_4_lut.init = 16'hcfc8;
    LUT4 i31985_2_lut_rep_926_3_lut (.A(n46143), .B(n46852), .C(n46155), 
         .Z(n46047)) /* synthesis lut_function=(A (B (C))+!A !(B+!(C))) */ ;
    defparam i31985_2_lut_rep_926_3_lut.init = 16'h9090;
    LUT4 i7335_2_lut_rep_991_4_lut_4_lut_4_lut (.A(n46125), .B(n93), .C(n46126), 
         .D(n124), .Z(n46112)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))+!B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i7335_2_lut_rep_991_4_lut_4_lut_4_lut.init = 16'h7662;
    LUT4 mux_86_i6_3_lut_rep_748_4_lut_4_lut (.A(n46003), .B(n45924), .C(n15), 
         .D(n45874), .Z(n45869)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_86_i6_3_lut_rep_748_4_lut_4_lut.init = 16'hc2c0;
    LUT4 i2_3_lut_adj_173 (.A(n45841), .B(n866[4]), .C(n45859), .Z(n41371)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i2_3_lut_adj_173.init = 16'h9696;
    LUT4 i2_4_lut_adj_174 (.A(n45861), .B(n754[2]), .C(n22446), .D(n21583), 
         .Z(n43695)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B !(D))) */ ;
    defparam i2_4_lut_adj_174.init = 16'h936c;
    LUT4 i1_2_lut_rep_795_4_lut (.A(n45925), .B(n73_adj_336), .C(n45926), 
         .D(n22673), .Z(n45916)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A (D)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_rep_795_4_lut.init = 16'hff08;
    LUT4 i4188_4_lut_4_lut (.A(n1429[1]), .B(n45796), .C(n580[2]), .D(n23030), 
         .Z(n6_adj_441)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !((D)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i4188_4_lut_4_lut.init = 16'h80ee;
    LUT4 i1_2_lut_rep_988_3_lut_3_lut_4_lut (.A(n46870), .B(n46127), .C(n29_adj_353), 
         .D(n46179), .Z(n46109)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_2_lut_rep_988_3_lut_3_lut_4_lut.init = 16'h0e00;
    LUT4 i37045_2_lut_rep_796_4_lut (.A(n15), .B(n46003), .C(n45924), 
         .D(n37_adj_301), .Z(n45917)) /* synthesis lut_function=(!(A ((D)+!B)+!A (((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i37045_2_lut_rep_796_4_lut.init = 16'h00c8;
    LUT4 i5787_4_lut_4_lut (.A(n1051[1]), .B(n1051[5]), .C(n1051[0]), 
         .D(n475[0]), .Z(n4_adj_370)) /* synthesis lut_function=(A ((C (D))+!B)+!A !(B+!(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5787_4_lut_4_lut.init = 16'hb332;
    LUT4 mux_47_i4_3_lut_rep_854_4_lut (.A(n46870), .B(n46127), .C(n45985), 
         .D(n46849), .Z(n45975)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam mux_47_i4_3_lut_rep_854_4_lut.init = 16'he0f1;
    LUT4 i6226_1_lut_3_lut_4_lut (.A(n46870), .B(n46127), .C(n45985), 
         .D(n46849), .Z(n8_adj_331)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i6226_1_lut_3_lut_4_lut.init = 16'h1f0e;
    CCU2D add_551_7 (.A0(VCC_net), .B0(n46016), .C0(n45777), .D0(n8965), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40491), 
          .S0(n2319[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_551_7.INIT0 = 16'ha956;
    defparam add_551_7.INIT1 = 16'h0000;
    defparam add_551_7.INJECT1_0 = "NO";
    defparam add_551_7.INJECT1_1 = "NO";
    LUT4 i17147_2_lut_rep_994_3_lut_4_lut (.A(n46128), .B(n89_adj_320), 
         .C(n89_adj_303), .D(n46145), .Z(n46115)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i17147_2_lut_rep_994_3_lut_4_lut.init = 16'h0200;
    CCU2D add_551_5 (.A0(n4445[2]), .B0(n45777), .C0(n825[7]), .D0(n46033), 
          .A1(n23068), .B1(n46033), .C1(n825[7]), .D1(n45777), .CIN(n40490), 
          .COUT(n40491), .S0(n2319[3]), .S1(n2319[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_551_5.INIT0 = 16'h5555;
    defparam add_551_5.INIT1 = 16'haaaa;
    defparam add_551_5.INJECT1_0 = "NO";
    defparam add_551_5.INJECT1_1 = "NO";
    LUT4 i14943_2_lut_4_lut (.A(n15), .B(n46003), .C(n45924), .D(n46077), 
         .Z(n4_adj_417)) /* synthesis lut_function=(!(A ((D)+!B)+!A (((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i14943_2_lut_4_lut.init = 16'h00c8;
    LUT4 i2_2_lut_rep_747_4_lut_4_lut (.A(n15), .B(n46003), .C(n45924), 
         .D(n45872), .Z(n45868)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B (C (D)+!C !(D))+!B !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i2_2_lut_rep_747_4_lut_4_lut.init = 16'hc297;
    LUT4 i63_else_4_lut_adj_175 (.A(akku_o_c_0), .B(n46189), .C(n117_adj_323), 
         .D(n122_adj_437), .Z(n46293)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i63_else_4_lut_adj_175.init = 16'h0001;
    LUT4 n334_bdd_2_lut_4_lut (.A(n45929), .B(n45940), .C(n37_adj_340), 
         .D(n46003), .Z(n45619)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (B+(C+(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam n334_bdd_2_lut_4_lut.init = 16'h00a3;
    LUT4 i2753_2_lut_rep_799_4_lut (.A(n45929), .B(n45940), .C(n37_adj_340), 
         .D(n46003), .Z(n45920)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (D)+!B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i2753_2_lut_rep_799_4_lut.init = 16'h5c00;
    CCU2D add_551_3 (.A0(n45781), .B0(n46033), .C0(n825[7]), .D0(n45777), 
          .A1(n8965), .B1(n8_adj_442), .C1(n23051), .D1(n46138), .CIN(n40489), 
          .COUT(n40490), .S0(n2319[1]), .S1(n2319[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_551_3.INIT0 = 16'haaaa;
    defparam add_551_3.INIT1 = 16'he111;
    defparam add_551_3.INJECT1_0 = "NO";
    defparam add_551_3.INJECT1_1 = "NO";
    LUT4 i5717_4_lut_4_lut (.A(n1582[1]), .B(n1582[5]), .C(n1582[0]), 
         .D(n615[0]), .Z(n4_adj_374)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5717_4_lut_4_lut.init = 16'heaa8;
    LUT4 i14910_2_lut_4_lut (.A(n45929), .B(n45940), .C(n37_adj_340), 
         .D(n46003), .Z(n21418)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B (D)+!B ((D)+!C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i14910_2_lut_4_lut.init = 16'hffa3;
    LUT4 mux_100_i3_3_lut (.A(n820), .B(n45816), .C(n15_adj_316), .Z(n429[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_100_i3_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_adj_176 (.A(n43753), .B(n45861), .C(n43695), .Z(n820)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i2_3_lut_adj_176.init = 16'h9696;
    LUT4 i14913_2_lut_rep_800_4_lut (.A(n45929), .B(n45940), .C(n37_adj_340), 
         .D(n46003), .Z(n45921)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A !(B+(C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i14913_2_lut_rep_800_4_lut.init = 16'ha300;
    LUT4 i23736_3_lut_4_lut_4_lut (.A(data[5]), .B(akku_o_c_8), .C(data[6]), 
         .D(data[7]), .Z(states_2__N_76[0])) /* synthesis lut_function=(!(A (C+(D))+!A !(B ((D)+!C)+!B !(C)))) */ ;
    defparam i23736_3_lut_4_lut_4_lut.init = 16'h450f;
    CCU2D add_551_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n43655), .B1(n43668), .C1(n46870), .D1(n45762), .COUT(n40489), 
          .S1(n2319[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_551_1.INIT0 = 16'hF000;
    defparam add_551_1.INIT1 = 16'h01ff;
    defparam add_551_1.INJECT1_0 = "NO";
    defparam add_551_1.INJECT1_1 = "NO";
    LUT4 mux_86_i3_4_lut (.A(n7_adj_443), .B(n330[2]), .C(n15), .D(n45572), 
         .Z(n363[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_86_i3_4_lut.init = 16'hcac5;
    LUT4 i2_3_lut_rep_801_4_lut (.A(n45975), .B(n45932), .C(n73_adj_336), 
         .D(n45925), .Z(n45922)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+!(C (D)))) */ ;
    defparam i2_3_lut_rep_801_4_lut.init = 16'h9000;
    LUT4 i2_4_lut_adj_177 (.A(n45862), .B(n23447), .C(n541[4]), .D(n330[2]), 
         .Z(n7_adj_443)) /* synthesis lut_function=(A (B)+!A !(B ((D)+!C)+!B !((D)+!C))) */ ;
    defparam i2_4_lut_adj_177.init = 16'h99c9;
    LUT4 mux_202_i7_3_lut_rep_650_4_lut (.A(n45779), .B(n46157), .C(n43563), 
         .D(n45773), .Z(n45771)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_202_i7_3_lut_rep_650_4_lut.init = 16'h08f8;
    LUT4 div_28_i85_3_lut_rep_996_4_lut_3_lut_4_lut_4_lut (.A(n46136), .B(n46132), 
         .C(n16[7]), .D(n93), .Z(n46117)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(B (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_i85_3_lut_rep_996_4_lut_3_lut_4_lut_4_lut.init = 16'h4c22;
    LUT4 i31366_2_lut_3_lut_4_lut (.A(n45779), .B(n46157), .C(n23081), 
         .D(n46130), .Z(n6_adj_355)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i31366_2_lut_3_lut_4_lut.init = 16'h0f8f;
    LUT4 div_53_i153_3_lut_4_lut_4_lut (.A(n45932), .B(n45961), .C(n45931), 
         .D(n191_adj_326), .Z(n220)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !(C+(D)))) */ ;
    defparam div_53_i153_3_lut_4_lut_4_lut.init = 16'hccc9;
    LUT4 n587_bdd_3_lut_4_lut (.A(n45888), .B(n45828), .C(n1429[1]), .D(n580[2]), 
         .Z(n45546)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+!(D)))+!A (C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam n587_bdd_3_lut_4_lut.init = 16'h0780;
    LUT4 i1_2_lut_rep_995_3_lut_3_lut_4_lut_4_lut (.A(n46136), .B(n46132), 
         .C(n16[7]), .D(n93), .Z(n46116)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B (D)+!B !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_rep_995_3_lut_3_lut_4_lut_4_lut.init = 16'h914c;
    LUT4 mux_72_i2_4_lut (.A(n5_adj_444), .B(n21[1]), .C(n43592), .D(n6_adj_407), 
         .Z(n3[1])) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_72_i2_4_lut.init = 16'h5cac;
    CCU2D div_39_add_172_7 (.A0(n4_adj_446), .B0(n45999), .C0(n45983), 
          .D0(n191), .A1(n45998), .B1(n45999), .C1(n45969), .D1(n190), 
          .CIN(n40487), .S0(n18[7]), .S1(n18[8]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_add_172_7.INIT0 = 16'h0ff4;
    defparam div_39_add_172_7.INIT1 = 16'h0bf4;
    defparam div_39_add_172_7.INJECT1_0 = "NO";
    defparam div_39_add_172_7.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_178 (.A(n45873), .B(n21395), .C(n21[1]), .D(n4_adj_393), 
         .Z(n5_adj_444)) /* synthesis lut_function=(!(A (B+(C (D)))+!A !(B+(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_4_lut_adj_178.init = 16'h5666;
    LUT4 i1_2_lut_rep_759_4_lut (.A(n3[8]), .B(n45933), .C(n6383), .D(n43720), 
         .Z(n45880)) /* synthesis lut_function=(A (B (D)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_rep_759_4_lut.init = 16'he817;
    CCU2D div_39_add_172_5 (.A0(n45981), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n45998), .B1(n45999), .C1(n45988), .D1(n46005), .CIN(n40486), 
          .COUT(n40487), .S0(n18[5]), .S1(n18[6]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_add_172_5.INIT0 = 16'h5555;
    defparam div_39_add_172_5.INIT1 = 16'h0bf4;
    defparam div_39_add_172_5.INJECT1_0 = "NO";
    defparam div_39_add_172_5.INJECT1_1 = "NO";
    LUT4 i14897_4_lut (.A(n45882), .B(n45867), .C(n45894), .D(n21[2]), 
         .Z(n21395)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D))+!B (C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i14897_4_lut.init = 16'h701a;
    LUT4 mux_47_i2_3_lut_4_lut (.A(n45937), .B(n43353), .C(n46123), .D(n107), 
         .Z(n107_adj_346)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_47_i2_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_65_i2_3_lut (.A(n40960), .B(n45902), .C(n37_adj_318), .Z(n21[1])) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_65_i2_3_lut.init = 16'h5c5c;
    LUT4 i2_2_lut_rep_613 (.A(n43673), .B(n7_adj_339), .Z(n45734)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i2_2_lut_rep_613.init = 16'h6666;
    LUT4 mux_195_i4_3_lut_4_lut (.A(n43673), .B(n7_adj_339), .C(n46157), 
         .D(n45743), .Z(n895[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam mux_195_i4_3_lut_4_lut.init = 16'hf909;
    LUT4 n45349_bdd_2_lut_3_lut (.A(n45348), .B(n270_adj_516[8]), .C(n270_adj_516[7]), 
         .Z(n45350)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam n45349_bdd_2_lut_3_lut.init = 16'hfefe;
    PFUMX i38764 (.BLUT(n46866), .ALUT(n46867), .C0(n43564), .Z(n43670));
    LUT4 i31361_2_lut_3_lut_4_lut (.A(n45779), .B(n46157), .C(n23081), 
         .D(n46130), .Z(n22564[2])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (C)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i31361_2_lut_3_lut_4_lut.init = 16'hf078;
    LUT4 i6_4_lut_adj_179 (.A(n9_adj_385), .B(n46170), .C(n46204), .D(n46205), 
         .Z(n15_adj_438)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam i6_4_lut_adj_179.init = 16'hfffe;
    CCU2D add_275_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n46261), .B1(n46264), .C1(n46229), .D1(n462[5]), .COUT(n40419), 
          .S1(n999[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_275_1.INIT0 = 16'hF000;
    defparam add_275_1.INIT1 = 16'h01ff;
    defparam add_275_1.INJECT1_0 = "NO";
    defparam add_275_1.INJECT1_1 = "NO";
    LUT4 i4_4_lut_adj_180 (.A(n7_adj_424), .B(n22867), .C(n45566), .D(n6_adj_414), 
         .Z(n40960)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i4_4_lut_adj_180.init = 16'h6996;
    PFUMX i38433 (.BLUT(n46287), .ALUT(n46288), .C0(n118_adj_307), .Z(n51_adj_344));
    CCU2D div_39_add_172_3 (.A0(n45998), .B0(n45999), .C0(n8_adj_451), 
          .D0(n46008), .A1(n45999), .B1(n46006), .C1(n45995), .D1(n45998), 
          .CIN(n40485), .COUT(n40486), .S0(n18[3]), .S1(n18[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_add_172_3.INIT0 = 16'h0b4f;
    defparam div_39_add_172_3.INIT1 = 16'hf072;
    defparam div_39_add_172_3.INJECT1_0 = "NO";
    defparam div_39_add_172_3.INJECT1_1 = "NO";
    LUT4 i5_4_lut_adj_181 (.A(n254), .B(n7_adj_452), .C(n250), .D(n8_adj_434), 
         .Z(n208[1])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i5_4_lut_adj_181.init = 16'hfffe;
    LUT4 i1_4_lut_adj_182 (.A(n255), .B(n251), .C(n107_adj_346), .D(n256), 
         .Z(n7_adj_452)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_182.init = 16'heccc;
    LUT4 i71_then_4_lut (.A(oprand[1]), .B(oprand[0]), .C(oprand[3]), 
         .D(oprand[2]), .Z(n46297)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i71_then_4_lut.init = 16'h0080;
    LUT4 i5_4_lut_adj_183 (.A(n254_adj_453), .B(n46382), .C(n251_adj_454), 
         .D(n8_adj_455), .Z(n146[1])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i5_4_lut_adj_183.init = 16'hfffe;
    LUT4 i1_2_lut_rep_1001_3_lut_4_lut (.A(n46870), .B(n43341), .C(n46145), 
         .D(n89_adj_320), .Z(n46122)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_2_lut_rep_1001_3_lut_4_lut.init = 16'h00e0;
    CCU2D div_39_add_172_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n46264), .B1(n46266), .C1(n112[2]), .D1(n112[4]), 
          .COUT(n40485), .S1(n18[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_add_172_1.INIT0 = 16'hF000;
    defparam div_39_add_172_1.INIT1 = 16'h0e1f;
    defparam div_39_add_172_1.INJECT1_0 = "NO";
    defparam div_39_add_172_1.INJECT1_1 = "NO";
    LUT4 mux_125_i4_3_lut_4_lut (.A(n46870), .B(n43341), .C(n45806), .D(n45804), 
         .Z(n545[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam mux_125_i4_3_lut_4_lut.init = 16'he0f1;
    LUT4 i15107_3_lut_rep_674_4_lut (.A(n45888), .B(n45828), .C(n580[2]), 
         .D(n1429[1]), .Z(n45795)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i15107_3_lut_rep_674_4_lut.init = 16'hf700;
    LUT4 i2_4_lut_adj_184 (.A(n45989), .B(n250_adj_456), .C(n18[6]), .D(n45951), 
         .Z(n8_adj_455)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;
    defparam i2_4_lut_adj_184.init = 16'hfcee;
    LUT4 akku_o_c_1_bdd_4_lut_38602 (.A(akku_o_c_1), .B(akku_o_c_3), .C(akku_o_c_2), 
         .D(akku_o_c_4), .Z(n46589)) /* synthesis lut_function=(A (B (C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D)))) */ ;
    defparam akku_o_c_1_bdd_4_lut_38602.init = 16'h9499;
    LUT4 mux_29_i2_3_lut (.A(n17[1]), .B(n248), .C(n7), .Z(n112[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_29_i2_3_lut.init = 16'hcaca;
    CCU2D add_502_7 (.A0(n2085[4]), .B0(n2085[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40484), 
          .S0(n2098[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_502_7.INIT0 = 16'h5999;
    defparam add_502_7.INIT1 = 16'h0000;
    defparam add_502_7.INJECT1_0 = "NO";
    defparam add_502_7.INJECT1_1 = "NO";
    CCU2D add_502_5 (.A0(n2085[2]), .B0(n2085[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2085[3]), .B1(n2085[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40483), .COUT(n40484), .S0(n2098[3]), .S1(n2098[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_502_5.INIT0 = 16'h5666;
    defparam add_502_5.INIT1 = 16'h5666;
    defparam add_502_5.INJECT1_0 = "NO";
    defparam add_502_5.INJECT1_1 = "NO";
    CCU2D add_502_3 (.A0(n2085[0]), .B0(n2085[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2085[1]), .B1(n2085[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40482), .COUT(n40483), .S0(n2098[1]), .S1(n2098[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_502_3.INIT0 = 16'h5999;
    defparam add_502_3.INIT1 = 16'h5999;
    defparam add_502_3.INJECT1_0 = "NO";
    defparam add_502_3.INJECT1_1 = "NO";
    LUT4 i6_4_lut_adj_185 (.A(n243), .B(n12_adj_457), .C(n30876), .D(n244), 
         .Z(n17[1])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut_adj_185.init = 16'hfffe;
    PFUMX i38378 (.BLUT(n45634), .ALUT(n45633), .C0(n6_adj_398), .Z(n45635));
    FD1P3AX pc_i0_i0 (.D(pc_5__N_35[0]), .SP(clk_c_enable_26), .CK(clk_c), 
            .Q(pc[0])) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam pc_i0_i0.GSR = "ENABLED";
    LUT4 mux_139_i5_3_lut_4_lut (.A(n45888), .B(n45828), .C(n46145), .D(n1416[1]), 
         .Z(n615[4])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_139_i5_3_lut_4_lut.init = 16'hf808;
    LUT4 i2179_4_lut_4_lut_4_lut (.A(n1[1]), .B(n22855), .C(n45939), .D(n23515), 
         .Z(n8_adj_400)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (B (C (D))+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2179_4_lut_4_lut_4_lut.init = 16'hfb20;
    LUT4 i5_4_lut_adj_186 (.A(n246_adj_458), .B(n242_adj_459), .C(n245), 
         .D(n241), .Z(n12_adj_457)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i5_4_lut_adj_186.init = 16'hfffe;
    LUT4 i2_3_lut_rep_808_4_lut (.A(n4201[1]), .B(n45935), .C(n6383), 
         .D(n3[8]), .Z(n45929)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C (D)))+!A (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_rep_808_4_lut.init = 16'h077f;
    CCU2D div_46_add_193_7 (.A0(n22712), .B0(n45965), .C0(n45949), .D0(n221_adj_435), 
          .A1(n22712), .B1(n45965), .C1(n45941), .D1(n220_adj_405), 
          .CIN(n40417), .S0(n270_adj_516[7]), .S1(n270_adj_516[8]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_46_add_193_7.INIT0 = 16'h0bf4;
    defparam div_46_add_193_7.INIT1 = 16'h0bf4;
    defparam div_46_add_193_7.INJECT1_0 = "NO";
    defparam div_46_add_193_7.INJECT1_1 = "NO";
    LUT4 i37134_3_lut_4_lut (.A(n46157), .B(n45), .C(n825[7]), .D(n46033), 
         .Z(n23081)) /* synthesis lut_function=(!((B+(C (D)+!C !(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i37134_3_lut_4_lut.init = 16'h0220;
    LUT4 i37246_3_lut_4_lut (.A(n46157), .B(n45), .C(n825[7]), .D(n46033), 
         .Z(n43991)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i37246_3_lut_4_lut.init = 16'h2220;
    CCU2D add_502_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(oprand[4]), .B1(oprand[3]), .C1(n5_adj_460), .D1(n720[1]), 
          .COUT(n40482), .S1(n2098[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_502_1.INIT0 = 16'hF000;
    defparam add_502_1.INIT1 = 16'h09ff;
    defparam add_502_1.INJECT1_0 = "NO";
    defparam add_502_1.INJECT1_1 = "NO";
    CCU2D add_500_7 (.A0(n2072[4]), .B0(n2072[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40481), 
          .S0(n2085[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_500_7.INIT0 = 16'h5999;
    defparam add_500_7.INIT1 = 16'h0000;
    defparam add_500_7.INJECT1_0 = "NO";
    defparam add_500_7.INJECT1_1 = "NO";
    LUT4 i4_4_lut_adj_187 (.A(n250_adj_461), .B(n251_adj_429), .C(n254_adj_430), 
         .D(n6_adj_462), .Z(n43353)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i4_4_lut_adj_187.init = 16'hfffe;
    CCU2D div_46_add_193_5 (.A0(n45950), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n45965), .B1(n45972), .C1(n22[6]), .D1(n22712), .CIN(n40416), 
          .COUT(n40417), .S0(n270_adj_516[5]), .S1(n270_adj_516[6]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_46_add_193_5.INIT0 = 16'h5555;
    defparam div_46_add_193_5.INIT1 = 16'h0f8d;
    defparam div_46_add_193_5.INJECT1_0 = "NO";
    defparam div_46_add_193_5.INJECT1_1 = "NO";
    CCU2D add_500_5 (.A0(n2072[2]), .B0(n2072[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2072[3]), .B1(n2072[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40480), .COUT(n40481), .S0(n2085[3]), .S1(n2085[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_500_5.INIT0 = 16'h5666;
    defparam add_500_5.INIT1 = 16'h5666;
    defparam add_500_5.INJECT1_0 = "NO";
    defparam add_500_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_897_3_lut_4_lut (.A(n46157), .B(n45), .C(n43563), 
         .D(n825[7]), .Z(n46018)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_897_3_lut_4_lut.init = 16'h0200;
    LUT4 mux_125_i3_3_lut_4_lut (.A(n45804), .B(n45800), .C(n46128), .D(n45803), 
         .Z(n545[2])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_125_i3_3_lut_4_lut.init = 16'hf606;
    CCU2D add_500_3 (.A0(n2072[0]), .B0(n2072[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2072[1]), .B1(n2072[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40479), .COUT(n40480), .S0(n2085[1]), .S1(n2085[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_500_3.INIT0 = 16'h5999;
    defparam add_500_3.INIT1 = 16'h5999;
    defparam add_500_3.INJECT1_0 = "NO";
    defparam add_500_3.INJECT1_1 = "NO";
    LUT4 i31356_2_lut_rep_655_3_lut_4_lut_4_lut (.A(n46157), .B(n45), .C(n825[7]), 
         .D(n45781), .Z(n45776)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i31356_2_lut_rep_655_3_lut_4_lut_4_lut.init = 16'h0200;
    LUT4 i24157_4_lut (.A(oprand[4]), .B(akku_o_c_4), .C(n46230), .D(n46229), 
         .Z(n3622)) /* synthesis lut_function=(A (B+(D))+!A (B (C)+!B (C (D)))) */ ;
    defparam i24157_4_lut.init = 16'hfac8;
    LUT4 i2241_2_lut_rep_915_3_lut_4_lut (.A(n46179), .B(n46064), .C(n23063), 
         .D(n46085), .Z(n46036)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i2241_2_lut_rep_915_3_lut_4_lut.init = 16'h0008;
    LUT4 i24252_2_lut_3_lut (.A(n43673), .B(n7_adj_339), .C(n23079), .Z(n30979)) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;
    defparam i24252_2_lut_3_lut.init = 16'hf6f6;
    CCU2D div_46_add_193_3 (.A0(n22712), .B0(n45971), .C0(n8_adj_464), 
          .D0(n45985), .A1(n254_adj_430), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n40415), .COUT(n40416), .S0(n270_adj_516[3]), 
          .S1(n270_adj_516[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_46_add_193_3.INIT0 = 16'hf4a0;
    defparam div_46_add_193_3.INIT1 = 16'h5555;
    defparam div_46_add_193_3.INJECT1_0 = "NO";
    defparam div_46_add_193_3.INJECT1_1 = "NO";
    LUT4 i2_3_lut_adj_188 (.A(n8_adj_465), .B(n45844), .C(n640[2]), .Z(n43732)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i2_3_lut_adj_188.init = 16'h9696;
    LUT4 i1_2_lut_4_lut_adj_189 (.A(n1416[1]), .B(n45827), .C(n45799), 
         .D(n45830), .Z(n23659)) /* synthesis lut_function=(A (B (C (D))+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_4_lut_adj_189.init = 16'ha200;
    LUT4 i1290_3_lut_rep_1012 (.A(states[0]), .B(\states[1] ), .C(n4_adj_440), 
         .Z(n46133)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(22[15:21])
    defparam i1290_3_lut_rep_1012.init = 16'h6262;
    CCU2D add_500_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(oprand[4]), .B1(oprand[3]), .C1(n5_adj_460), .D1(n45763), 
          .COUT(n40479), .S1(n2085[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_500_1.INIT0 = 16'hF000;
    defparam add_500_1.INIT1 = 16'h09ff;
    defparam add_500_1.INJECT1_0 = "NO";
    defparam add_500_1.INJECT1_1 = "NO";
    LUT4 akku_o_c_1_bdd_4_lut_38603 (.A(akku_o_c_1), .B(akku_o_c_3), .C(akku_o_c_2), 
         .D(akku_o_c_4), .Z(n106_adj_312)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;
    defparam akku_o_c_1_bdd_4_lut_38603.init = 16'h0db0;
    LUT4 i23839_2_lut_rep_928_3_lut (.A(n46143), .B(n46852), .C(n46155), 
         .Z(n46049)) /* synthesis lut_function=(!(A (B (C))+!A !(B+!(C)))) */ ;
    defparam i23839_2_lut_rep_928_3_lut.init = 16'h6f6f;
    LUT4 mux_132_i4_3_lut_rep_678 (.A(n1298[5]), .B(n545[3]), .C(n89_adj_320), 
         .Z(n45799)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_132_i4_3_lut_rep_678.init = 16'h5c5c;
    LUT4 i1_4_lut_adj_190 (.A(n45812), .B(n41282), .C(n45809), .D(n6_adj_466), 
         .Z(n43738)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+!(D)))+!A !(B ((D)+!C)+!B !(C+!(D))))) */ ;
    defparam i1_4_lut_adj_190.init = 16'h65a6;
    LUT4 i4133_2_lut_4_lut (.A(n1298[5]), .B(n545[3]), .C(n89_adj_320), 
         .D(n45827), .Z(n1429[1])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(B (D)+!B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i4133_2_lut_4_lut.init = 16'ha35c;
    LUT4 n863_bdd_3_lut_rep_635_4_lut (.A(n45781), .B(n45), .C(n45758), 
         .D(n860[5]), .Z(n45756)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam n863_bdd_3_lut_rep_635_4_lut.init = 16'h2000;
    LUT4 i2582_3_lut_4_lut_4_lut_4_lut_4_lut (.A(n46014), .B(n45940), .C(n3[4]), 
         .D(n45929), .Z(n6_adj_416)) /* synthesis lut_function=(!(A (B)+!A !(B (C+!(D))+!B !((D)+!C)))) */ ;
    defparam i2582_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h6276;
    LUT4 i1_2_lut_rep_676_4_lut (.A(n45890), .B(n6_adj_402), .C(n8_adj_401), 
         .D(n45804), .Z(n45797)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i1_2_lut_rep_676_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_992_3_lut_4_lut_4_lut (.A(n16[7]), .B(n16[8]), .C(n46870), 
         .D(n7), .Z(n46113)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !((C+!(D))+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_992_3_lut_4_lut_4_lut.init = 16'hac80;
    LUT4 i2_4_lut_adj_191 (.A(n21590), .B(n22969), .C(n23490), .D(n45832), 
         .Z(n43753)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B (C (D))+!B !(C (D)))) */ ;
    defparam i2_4_lut_adj_191.init = 16'h9666;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n46014), .B(n45940), .C(n3[4]), 
         .D(n45929), .Z(n22902)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !((D)+!C))+!A !(B (C+!(D))+!B !((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h6a56;
    LUT4 akku_o_c_1_bdd_4_lut_38742 (.A(akku_o_c_1), .B(akku_o_c_3), .C(akku_o_c_2), 
         .D(akku_o_c_4), .Z(n46151)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+!(D)))+!A !(B ((D)+!C)+!B (C+!(D)))) */ ;
    defparam akku_o_c_1_bdd_4_lut_38742.init = 16'h83c8;
    LUT4 i1_2_lut_4_lut_adj_192 (.A(n1169[2]), .B(n45804), .C(n45802), 
         .D(n43678), .Z(n4_adj_467)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_4_lut_adj_192.init = 16'h57a8;
    LUT4 mux_132_i2_3_lut (.A(n1324[5]), .B(n545[1]), .C(n89_adj_320), 
         .Z(n580[1])) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_132_i2_3_lut.init = 16'h5c5c;
    LUT4 mux_125_i2_4_lut (.A(n45800), .B(n510[1]), .C(n46128), .D(n4_adj_467), 
         .Z(n545[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_125_i2_4_lut.init = 16'hcac5;
    LUT4 mux_153_i5_3_lut_4_lut (.A(n46144), .B(n46870), .C(n45794), .D(n1687[5]), 
         .Z(n685[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam mux_153_i5_3_lut_4_lut.init = 16'he0f1;
    LUT4 i37240_2_lut_rep_701_3_lut_4_lut (.A(n46144), .B(n46870), .C(n89_adj_303), 
         .D(n45829), .Z(n45822)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i37240_2_lut_rep_701_3_lut_4_lut.init = 16'h0e00;
    LUT4 mux_153_i3_3_lut_4_lut (.A(n46144), .B(n46870), .C(n650[2]), 
         .D(n45774), .Z(n685[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam mux_153_i3_3_lut_4_lut.init = 16'he0f1;
    LUT4 i1_4_lut_adj_193 (.A(n22998), .B(n40801), .C(n7458), .D(n7_adj_468), 
         .Z(n43678)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A !(B (C+!(D))+!B (C)))) */ ;
    defparam i1_4_lut_adj_193.init = 16'h5a56;
    LUT4 i3347_4_lut (.A(n45797), .B(n45801), .C(n22887), .D(n510[1]), 
         .Z(n7458)) /* synthesis lut_function=(!((B+!((D)+!C))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3347_4_lut.init = 16'h2202;
    LUT4 i3872_4_lut_4_lut (.A(n1169[2]), .B(n45804), .C(n45802), .D(n22998), 
         .Z(n8_adj_401)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A (B+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3872_4_lut_4_lut.init = 16'h20bb;
    LUT4 i2_2_lut_3_lut_4_lut_adj_194 (.A(n1169[2]), .B(n45804), .C(n45802), 
         .D(n45800), .Z(n7_adj_469)) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (D)+!B !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_2_lut_3_lut_4_lut_adj_194.init = 16'h9b64;
    LUT4 mux_118_i2_3_lut (.A(n1051[5]), .B(n475[1]), .C(n45_adj_356), 
         .Z(n510[1])) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_118_i2_3_lut.init = 16'h5c5c;
    LUT4 i71_else_4_lut (.A(oprand[1]), .B(oprand[0]), .C(oprand[3]), 
         .D(oprand[2]), .Z(n46296)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i71_else_4_lut.init = 16'h0001;
    LUT4 i37088_2_lut_rep_660_3_lut_4_lut (.A(n46870), .B(n46146), .C(n43564), 
         .D(n755[6]), .Z(n45781)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i37088_2_lut_rep_660_3_lut_4_lut.init = 16'h0e00;
    LUT4 i4_4_lut_adj_195 (.A(n41371), .B(n43741), .C(n43738), .D(n6_adj_470), 
         .Z(n910[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i4_4_lut_adj_195.init = 16'h6996;
    LUT4 i1_2_lut_3_lut_4_lut_adj_196 (.A(n45805), .B(n45804), .C(n45803), 
         .D(n45800), .Z(n7_adj_468)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B (D)+!B !((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_196.init = 16'h4412;
    LUT4 mux_181_i5_3_lut_4_lut (.A(n46870), .B(n46146), .C(n790[4]), 
         .D(n2203[5]), .Z(n825[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam mux_181_i5_3_lut_4_lut.init = 16'he0f1;
    LUT4 mux_100_i2_4_lut (.A(n7_adj_471), .B(n396[1]), .C(n15_adj_316), 
         .D(n8_adj_472), .Z(n429[1])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_100_i2_4_lut.init = 16'hc5ca;
    LUT4 i2_4_lut_adj_197 (.A(n776[2]), .B(n41143), .C(n40708), .D(n30785), 
         .Z(n7_adj_471)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C (D))+!B !((D)+!C)))) */ ;
    defparam i2_4_lut_adj_197.init = 16'h6a9a;
    LUT4 i3_4_lut_adj_198 (.A(n43753), .B(n41286), .C(n23490), .D(n45814), 
         .Z(n8_adj_472)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B (C (D)+!C !(D))+!B !(C))) */ ;
    defparam i3_4_lut_adj_198.init = 16'h965a;
    LUT4 i2_4_lut_adj_199 (.A(n45816), .B(n396[1]), .C(n41286), .D(n820), 
         .Z(n40708)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_4_lut_adj_199.init = 16'hffde;
    CCU2D add_498_7 (.A0(n2059[4]), .B0(n2059[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40478), 
          .S0(n2072[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_498_7.INIT0 = 16'h5999;
    defparam add_498_7.INIT1 = 16'h0000;
    defparam add_498_7.INJECT1_0 = "NO";
    defparam add_498_7.INJECT1_1 = "NO";
    LUT4 i3_4_lut_4_lut_adj_200 (.A(n46150), .B(n46880), .C(n31204), .D(n46339), 
         .Z(n7)) /* synthesis lut_function=(A (B+(C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i3_4_lut_4_lut_adj_200.init = 16'hffbd;
    LUT4 i1_4_lut_adj_201 (.A(n6_adj_466), .B(n41354), .C(n45807), .D(n6_adj_373), 
         .Z(n43741)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B (C+!(D))+!B !((D)+!C))) */ ;
    defparam i1_4_lut_adj_201.init = 16'h95a9;
    LUT4 i4472_4_lut_4_lut (.A(n45784), .B(n45782), .C(n650[2]), .D(n45785), 
         .Z(n6_adj_422)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i4472_4_lut_4_lut.init = 16'hee80;
    LUT4 i23734_4_lut (.A(n46282), .B(n46138), .C(n755[0]), .D(n43564), 
         .Z(n825[0])) /* synthesis lut_function=(A (B (C+(D)))+!A !(((D)+!C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i23734_4_lut.init = 16'h88c0;
    CCU2D add_498_5 (.A0(n2059[2]), .B0(n2059[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2059[3]), .B1(n2059[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40477), .COUT(n40478), .S0(n2072[3]), .S1(n2072[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_498_5.INIT0 = 16'h5666;
    defparam add_498_5.INIT1 = 16'h5666;
    defparam add_498_5.INJECT1_0 = "NO";
    defparam add_498_5.INJECT1_1 = "NO";
    CCU2D div_46_add_193_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n45957), .B1(n45958), .C1(n11), .D1(n45974), 
          .COUT(n40415), .S1(n270_adj_516[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_46_add_193_1.INIT0 = 16'hF000;
    defparam div_46_add_193_1.INIT1 = 16'h01f1;
    defparam div_46_add_193_1.INJECT1_0 = "NO";
    defparam div_46_add_193_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_202 (.A(n45825), .B(n43727), .C(n45819), .D(n6_adj_378), 
         .Z(n43765)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+!(D)))+!A !(B ((D)+!C)+!B !(C+!(D))))) */ ;
    defparam i1_4_lut_adj_202.init = 16'h65a6;
    LUT4 i2_3_lut_4_lut_adj_203 (.A(n45805), .B(n45803), .C(n1169[2]), 
         .D(n45804), .Z(n40801)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C (D)+!C !(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_4_lut_adj_203.init = 16'h0f1e;
    CCU2D add_498_3 (.A0(n2059[0]), .B0(n2059[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2059[1]), .B1(n2059[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40476), .COUT(n40477), .S0(n2072[1]), .S1(n2072[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_498_3.INIT0 = 16'h5999;
    defparam add_498_3.INIT1 = 16'h5999;
    defparam add_498_3.INJECT1_0 = "NO";
    defparam add_498_3.INJECT1_1 = "NO";
    LUT4 akku_o_c_0_bdd_3_lut (.A(akku_o_c_0), .B(akku_o_c_4), .C(akku_o_c_3), 
         .Z(n45374)) /* synthesis lut_function=(A (B (C))+!A !(B+(C))) */ ;
    defparam akku_o_c_0_bdd_3_lut.init = 16'h8181;
    LUT4 mux_118_i3_3_lut_rep_682 (.A(n1038[5]), .B(n475[2]), .C(n45_adj_356), 
         .Z(n45803)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_118_i3_3_lut_rep_682.init = 16'h5c5c;
    LUT4 n43564_bdd_4_lut_4_lut (.A(n755[6]), .B(n43564), .C(n755[5]), 
         .D(n46040), .Z(n2203[5])) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam n43564_bdd_4_lut_4_lut.init = 16'hdfff;
    LUT4 i2_3_lut_adj_204 (.A(n363[2]), .B(n41291), .C(n45848), .Z(n41388)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i2_3_lut_adj_204.init = 16'h9696;
    PFUMX i38373 (.BLUT(n45627), .ALUT(n45626), .C0(n45759), .Z(n6_adj_398));
    LUT4 i1_2_lut_4_lut_adj_205 (.A(n1038[5]), .B(n475[2]), .C(n45_adj_356), 
         .D(n45804), .Z(n22887)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(B (D)+!B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_4_lut_adj_205.init = 16'ha35c;
    LUT4 i37194_3_lut_4_lut (.A(akku_o_c_1), .B(n46151), .C(n106_adj_312), 
         .D(n110_adj_311), .Z(n32)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;
    defparam i37194_3_lut_4_lut.init = 16'h0009;
    LUT4 i3858_2_lut_rep_681_4_lut (.A(n1038[5]), .B(n475[2]), .C(n45_adj_356), 
         .D(n45805), .Z(n45802)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A (B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i3858_2_lut_rep_681_4_lut.init = 16'hff5c;
    CCU2D add_498_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n43701), .B1(n7_adj_397), .C1(n19), .D1(n46847), .COUT(n40476), 
          .S1(n2072[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_498_1.INIT0 = 16'hF000;
    defparam add_498_1.INIT1 = 16'h06f6;
    defparam add_498_1.INJECT1_0 = "NO";
    defparam add_498_1.INJECT1_1 = "NO";
    CCU2D add_496_7 (.A0(n2046[4]), .B0(n2046[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40475), 
          .S0(n2059[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_496_7.INIT0 = 16'h5999;
    defparam add_496_7.INIT1 = 16'h0000;
    defparam add_496_7.INJECT1_0 = "NO";
    defparam add_496_7.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_206 (.A(n46235), .B(n103), .C(n43606), .D(n46376), 
         .Z(n89_adj_303)) /* synthesis lut_function=(A (B (D))+!A !((C+!(D))+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_4_lut_adj_206.init = 16'h8c00;
    LUT4 i24147_2_lut_rep_883_3_lut_4_lut_4_lut (.A(n46155), .B(n217), .C(n22715), 
         .D(n46049), .Z(n46004)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C+!(D))))) */ ;
    defparam i24147_2_lut_rep_883_3_lut_4_lut_4_lut.init = 16'h4844;
    LUT4 i1_2_lut_rep_870_3_lut_4_lut_4_lut (.A(n46155), .B(n217), .C(n22716), 
         .D(n46029), .Z(n45991)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (C+!(D))+!B (C))) */ ;
    defparam i1_2_lut_rep_870_3_lut_4_lut_4_lut.init = 16'hf8f4;
    CCU2D add_496_5 (.A0(n2046[2]), .B0(n2046[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2046[3]), .B1(n2046[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40474), .COUT(n40475), .S0(n2059[3]), .S1(n2059[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_496_5.INIT0 = 16'h5666;
    defparam add_496_5.INIT1 = 16'h5666;
    defparam add_496_5.INJECT1_0 = "NO";
    defparam add_496_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_207 (.A(akku_o_c_4), .B(akku_o_c_3), .Z(n43606)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i1_2_lut_adj_207.init = 16'h2222;
    CCU2D add_496_3 (.A0(n2046[0]), .B0(n2046[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n2046[1]), .B1(n2046[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40473), .COUT(n40474), .S0(n2059[1]), .S1(n2059[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_496_3.INIT0 = 16'h5999;
    defparam add_496_3.INIT1 = 16'h5999;
    defparam add_496_3.INJECT1_0 = "NO";
    defparam add_496_3.INJECT1_1 = "NO";
    LUT4 i5065_2_lut_rep_656_3_lut_4_lut (.A(n46138), .B(n45783), .C(n2293[1]), 
         .D(n825[7]), .Z(n45777)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A !((D)+!C)) */ ;
    defparam i5065_2_lut_rep_656_3_lut_4_lut.init = 16'h80f0;
    LUT4 i5063_2_lut_3_lut_4_lut (.A(n46138), .B(n45783), .C(n2293[1]), 
         .D(n825[7]), .Z(n4445[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;
    defparam i5063_2_lut_3_lut_4_lut.init = 16'h780f;
    CCU2D div_39_add_193_9 (.A0(n45957), .B0(n45958), .C0(n18[7]), .D0(n221), 
          .A1(n45957), .B1(n45958), .C1(n18[8]), .D1(n45964), .CIN(n40413), 
          .S0(n270_adj_514[7]), .S1(n270_adj_514[8]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_add_193_9.INIT0 = 16'h0e1f;
    defparam div_39_add_193_9.INIT1 = 16'h0e1f;
    defparam div_39_add_193_9.INJECT1_0 = "NO";
    defparam div_39_add_193_9.INJECT1_1 = "NO";
    LUT4 div_53_i156_3_lut_3_lut_4_lut_4_lut (.A(n45946), .B(n41038), .C(n45953), 
         .D(n45945), .Z(n223)) /* synthesis lut_function=(A (B)+!A (B ((D)+!C)+!B !(C+(D)))) */ ;
    defparam div_53_i156_3_lut_3_lut_4_lut_4_lut.init = 16'hcc8d;
    LUT4 i1_2_lut_rep_900_3_lut_4_lut_3_lut (.A(n46155), .B(n22715), .C(n46057), 
         .Z(n46021)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;
    defparam i1_2_lut_rep_900_3_lut_4_lut_3_lut.init = 16'h6464;
    LUT4 i1_2_lut_rep_936_4_lut (.A(n16[4]), .B(n16[5]), .C(n46870), .D(n46852), 
         .Z(n46057)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_936_4_lut.init = 16'h53ac;
    LUT4 mux_54_i4_3_lut_3_lut_4_lut_4_lut (.A(n45946), .B(n29_adj_353), 
         .C(n45975), .D(n45945), .Z(n218[3])) /* synthesis lut_function=(A (B+(C))+!A (B (D)+!B (C))) */ ;
    defparam mux_54_i4_3_lut_3_lut_4_lut_4_lut.init = 16'hfcb8;
    LUT4 i1_2_lut_4_lut_adj_208 (.A(n6_adj_402), .B(n46051), .C(n45896), 
         .D(n43678), .Z(n43679)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (D)+!B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_4_lut_adj_208.init = 16'h8976;
    LUT4 i38138_2_lut_rep_1023 (.A(n44162), .B(n44765), .Z(n46144)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i38138_2_lut_rep_1023.init = 16'heeee;
    LUT4 i2165_4_lut_3_lut_rep_818 (.A(n22855), .B(n45947), .C(n45987), 
         .Z(n45939)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2165_4_lut_3_lut_rep_818.init = 16'h8e8e;
    CCU2D add_496_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n45760), .B1(n45765), .C1(n19), .D1(n45791), .COUT(n40473), 
          .S1(n2059[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_496_1.INIT0 = 16'hF000;
    defparam add_496_1.INIT1 = 16'h01f1;
    defparam add_496_1.INJECT1_0 = "NO";
    defparam add_496_1.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_209 (.A(n8_adj_476), .B(n22896), .C(n45821), .D(n45793), 
         .Z(n23779)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B ((D)+!C)+!B !((D)+!C))) */ ;
    defparam i2_4_lut_adj_209.init = 16'h9969;
    LUT4 i2172_3_lut_rep_807_3_lut_4_lut (.A(n22855), .B(n45947), .C(n45987), 
         .D(n1[1]), .Z(n45928)) /* synthesis lut_function=(A (B+((D)+!C))+!A !((C+!(D))+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2172_3_lut_rep_807_3_lut_4_lut.init = 16'hae8a;
    LUT4 i4444_4_lut (.A(n45793), .B(n1687[5]), .C(n45821), .D(n6_adj_376), 
         .Z(n8_adj_476)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !((D)+!C))+!A !(B (C (D))+!B (C+(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i4444_4_lut.init = 16'h7b12;
    CCU2D add_494_7 (.A0(VCC_net), .B0(n46026), .C0(n46040), .D0(n38250), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40472), 
          .S0(n2046[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_494_7.INIT0 = 16'ha955;
    defparam add_494_7.INIT1 = 16'h0000;
    defparam add_494_7.INJECT1_0 = "NO";
    defparam add_494_7.INJECT1_1 = "NO";
    LUT4 mux_139_i4_3_lut_4_lut (.A(n45481), .B(n46147), .C(n45799), .D(n45831), 
         .Z(n615[3])) /* synthesis lut_function=(A (C)+!A !(B (D)+!B !(C))) */ ;
    defparam mux_139_i4_3_lut_4_lut.init = 16'hb0f4;
    LUT4 i2_3_lut_rep_934_4_lut (.A(n45481), .B(n46147), .C(n46066), .D(n89_adj_320), 
         .Z(n46055)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B+((D)+!C)))) */ ;
    defparam i2_3_lut_rep_934_4_lut.init = 16'h00b0;
    LUT4 i1_2_lut_rep_1025 (.A(n43655), .B(n43668), .Z(n46146)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_2_lut_rep_1025.init = 16'heeee;
    LUT4 i2_3_lut_4_lut_adj_210 (.A(n22855), .B(n45947), .C(n45987), .D(n1[1]), 
         .Z(n41244)) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_4_lut_adj_210.init = 16'hdb24;
    LUT4 i1_2_lut_3_lut_4_lut_adj_211 (.A(n43655), .B(n43668), .C(n43564), 
         .D(n46870), .Z(n43581)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_2_lut_3_lut_4_lut_adj_211.init = 16'h0f0e;
    CCU2D add_494_5 (.A0(n45264), .B0(n755[6]), .C0(n46040), .D0(n46026), 
          .A1(n44022), .B1(n755[6]), .C1(n46040), .D1(n46026), .CIN(n40471), 
          .COUT(n40472), .S0(n2046[3]), .S1(n2046[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_494_5.INIT0 = 16'h5555;
    defparam add_494_5.INIT1 = 16'h5555;
    defparam add_494_5.INJECT1_0 = "NO";
    defparam add_494_5.INJECT1_1 = "NO";
    LUT4 i2_4_lut_else_4_lut_adj_212 (.A(n2098[5]), .B(n2098[4]), .C(n2098[2]), 
         .D(n4_adj_347), .Z(n46280)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B)) */ ;
    defparam i2_4_lut_else_4_lut_adj_212.init = 16'hccc6;
    LUT4 div_46_i174_3_lut_4_lut (.A(n221_adj_435), .B(n45949), .C(n45966), 
         .D(n220_adj_405), .Z(n250_adj_461)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_46_i174_3_lut_4_lut.init = 16'hfe01;
    LUT4 i24320_2_lut_3_lut_4_lut (.A(n46214), .B(n46160), .C(akku_o_c_0), 
         .D(akku_o_c_1), .Z(n31047)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i24320_2_lut_3_lut_4_lut.init = 16'hf1fe;
    CCU2D add_494_3 (.A0(n46015), .B0(n8_adj_477), .C0(n755[6]), .D0(GND_net), 
          .A1(n46015), .B1(n8_adj_477), .C1(n755[6]), .D1(n46040), .CIN(n40470), 
          .COUT(n40471), .S0(n2046[1]), .S1(n2046[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_494_3.INIT0 = 16'hee1e;
    defparam add_494_3.INIT1 = 16'he11e;
    defparam add_494_3.INJECT1_0 = "NO";
    defparam add_494_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_213 (.A(n46214), .B(n46160), .C(akku_o_c_0), 
         .D(akku_o_c_1), .Z(n41396)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i1_2_lut_3_lut_4_lut_adj_213.init = 16'h1ee1;
    LUT4 i15336_2_lut_4_lut_4_lut_4_lut (.A(n45952), .B(n45975), .C(n45926), 
         .D(n45932), .Z(n22035)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B (C+!(D))+!B (C)))) */ ;
    defparam i15336_2_lut_4_lut_4_lut_4_lut.init = 16'h0509;
    LUT4 i1_3_lut_rep_680_4_lut (.A(n45806), .B(n45891), .C(n45803), .D(n45804), 
         .Z(n45801)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_3_lut_rep_680_4_lut.init = 16'h9996;
    LUT4 i23985_2_lut_rep_816_4_lut (.A(n45951), .B(n45974), .C(n11), 
         .D(n45948), .Z(n45937)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i23985_2_lut_rep_816_4_lut.init = 16'h00ca;
    LUT4 i15073_3_lut_4_lut (.A(n1156[1]), .B(n45806), .C(n45891), .D(n1156[2]), 
         .Z(n6_adj_402)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i15073_3_lut_4_lut.init = 16'hef00;
    LUT4 i2_3_lut_4_lut_adj_214 (.A(n1156[1]), .B(n45806), .C(n1156[2]), 
         .D(n45891), .Z(n22998)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_4_lut_adj_214.init = 16'he1f0;
    LUT4 i24365_3_lut_4_lut (.A(n118_adj_307), .B(n46164), .C(n5), .D(n117_adj_305), 
         .Z(n122_adj_375)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i24365_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_118_i4_3_lut_rep_685 (.A(n1025[5]), .B(n475[3]), .C(n45_adj_356), 
         .Z(n45806)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_118_i4_3_lut_rep_685.init = 16'h5c5c;
    LUT4 i2_4_lut_adj_215 (.A(n45783), .B(n8_adj_342), .C(n45762), .D(n46364), 
         .Z(n23806)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i2_4_lut_adj_215.init = 16'h6996;
    LUT4 i3_2_lut_3_lut_4_lut (.A(n46166), .B(n46165), .C(n46167), .D(n46168), 
         .Z(n9_adj_478)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 oprand_2__bdd_4_lut (.A(n46882), .B(n46878), .C(n46873), .D(n46875), 
         .Z(n46790)) /* synthesis lut_function=(A (B (C (D))+!B !(C+!(D)))+!A !(B ((D)+!C)+!B (C+(D)))) */ ;
    defparam oprand_2__bdd_4_lut.init = 16'h8241;
    LUT4 i2_3_lut_adj_216 (.A(n45757), .B(n2203[5]), .C(n790[4]), .Z(n2216[2])) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_adj_216.init = 16'h1e1e;
    LUT4 i37196_3_lut_4_lut (.A(oprand[1]), .B(n46159), .C(n106), .D(n110), 
         .Z(n23)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A ((C+(D))+!B))) */ ;
    defparam i37196_3_lut_4_lut.init = 16'h0006;
    LUT4 i2_2_lut_rep_1168 (.A(\states[1] ), .B(states[0]), .C(n4_adj_440), 
         .Z(n46854)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam i2_2_lut_rep_1168.init = 16'h0202;
    LUT4 i3810_2_lut_rep_684_4_lut (.A(n1025[5]), .B(n475[3]), .C(n45_adj_356), 
         .D(n45891), .Z(n45805)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(B (D)+!B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i3810_2_lut_rep_684_4_lut.init = 16'ha35c;
    LUT4 i32049_2_lut_rep_810_3_lut_4_lut_4_lut_4_lut (.A(n45953), .B(n45975), 
         .C(n45954), .D(n45952), .Z(n45931)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;
    defparam i32049_2_lut_rep_810_3_lut_4_lut_4_lut_4_lut.init = 16'hf0f4;
    CCU2D add_494_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n46847), .B1(n45791), .C1(n19), .D1(n720[5]), .COUT(n40470), 
          .S1(n2046[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_494_1.INIT0 = 16'hF000;
    defparam add_494_1.INIT1 = 16'h0dff;
    defparam add_494_1.INJECT1_0 = "NO";
    defparam add_494_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_217 (.A(n45725), .B(n43706), .Z(n43708)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_adj_217.init = 16'h6666;
    LUT4 i32057_2_lut_rep_806_3_lut_4_lut_4_lut (.A(n45953), .B(n45954), 
         .C(n191_adj_326), .D(n45938), .Z(n45927)) /* synthesis lut_function=(A (B+(C))+!A (B+(C+(D)))) */ ;
    defparam i32057_2_lut_rep_806_3_lut_4_lut_4_lut.init = 16'hfdfc;
    LUT4 i15810_4_lut_4_lut (.A(\states[1] ), .B(states[0]), .C(n4_adj_440), 
         .D(akku_o_8__N_50[5]), .Z(n22537)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam i15810_4_lut_4_lut.init = 16'hfd00;
    LUT4 i2_3_lut_4_lut_adj_218 (.A(n429[2]), .B(n45807), .C(n429[1]), 
         .D(n23471), .Z(n41383)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_4_lut_adj_218.init = 16'h42bd;
    LUT4 mux_195_i5_3_lut_4_lut (.A(n46177), .B(n43349), .C(n45758), .D(n2476[5]), 
         .Z(n895[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam mux_195_i5_3_lut_4_lut.init = 16'he0f1;
    LUT4 i1_2_lut_rep_805_3_lut_4_lut_4_lut_4_lut_4_lut_4_lut (.A(n45953), 
         .B(n45946), .C(n45975), .D(n45952), .Z(n45926)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B (C)+!B !(C (D)))) */ ;
    defparam i1_2_lut_rep_805_3_lut_4_lut_4_lut_4_lut_4_lut_4_lut.init = 16'hc3d3;
    CCU2D div_39_add_193_7 (.A0(n45957), .B0(n45958), .C0(n18[5]), .D0(n45981), 
          .A1(n45957), .B1(n45958), .C1(n18[6]), .D1(n45989), .CIN(n40412), 
          .COUT(n40413), .S0(n270_adj_514[5]), .S1(n270_adj_514[6]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_add_193_7.INIT0 = 16'h0e1f;
    defparam div_39_add_193_7.INIT1 = 16'h0e1f;
    defparam div_39_add_193_7.INJECT1_0 = "NO";
    defparam div_39_add_193_7.INJECT1_1 = "NO";
    LUT4 i1301_2_lut_rep_1155 (.A(\states[1] ), .B(states[0]), .Z(n46276)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam i1301_2_lut_rep_1155.init = 16'h2222;
    LUT4 i2_4_lut_adj_219 (.A(n21806), .B(n2476[5]), .C(n30979), .D(n2476[3]), 
         .Z(n43712)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i2_4_lut_adj_219.init = 16'h9c63;
    LUT4 i15168_4_lut (.A(n2476[5]), .B(n21805), .C(n2476[2]), .D(n22479), 
         .Z(n21806)) /* synthesis lut_function=(!(A ((C (D)+!C !(D))+!B)+!A ((C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i15168_4_lut.init = 16'h0c84;
    LUT4 i1_2_lut_rep_1009_4_lut (.A(n46177), .B(n43349), .C(n825[7]), 
         .D(n45), .Z(n46130)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_2_lut_rep_1009_4_lut.init = 16'h00e0;
    LUT4 i5037_4_lut (.A(n45734), .B(n2489[1]), .C(n23079), .D(n860[1]), 
         .Z(n21805)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5037_4_lut.init = 16'h5f5d;
    LUT4 mux_181_i2_4_lut (.A(n43709), .B(n790[1]), .C(n46138), .D(n4_adj_351), 
         .Z(n825[1])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_181_i2_4_lut.init = 16'hc5ca;
    CCU2D div_39_add_193_5 (.A0(n45992), .B0(n46008), .C0(n18[3]), .D0(n45951), 
          .A1(n45963), .B1(n45957), .C1(n18[4]), .D1(n224), .CIN(n40411), 
          .COUT(n40412), .S0(n270_adj_514[3]), .S1(n270_adj_514[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_add_193_5.INIT0 = 16'hf099;
    defparam div_39_add_193_5.INIT1 = 16'h0e3f;
    defparam div_39_add_193_5.INJECT1_0 = "NO";
    defparam div_39_add_193_5.INJECT1_1 = "NO";
    CCU2D div_39_add_193_3 (.A0(n46264), .B0(n46266), .C0(n112[1]), .D0(n112[3]), 
          .A1(n45957), .B1(n45958), .C1(n18[2]), .D1(n45974), .CIN(n40410), 
          .COUT(n40411), .S0(n270_adj_514[1]), .S1(n270_adj_514[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_add_193_3.INIT0 = 16'hf1e0;
    defparam div_39_add_193_3.INIT1 = 16'h0e1f;
    defparam div_39_add_193_3.INJECT1_0 = "NO";
    defparam div_39_add_193_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_220 (.A(n46138), .B(n45783), .C(n860[5]), 
         .D(n45), .Z(n23070)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_220.init = 16'hf078;
    LUT4 oprand_4__bdd_4_lut_38535 (.A(n46873), .B(oprand[3]), .C(oprand[2]), 
         .D(oprand[1]), .Z(n9_adj_484)) /* synthesis lut_function=(!((B (C (D)))+!A)) */ ;
    defparam oprand_4__bdd_4_lut_38535.init = 16'h2aaa;
    LUT4 mux_174_i2_4_lut (.A(n2098[5]), .B(n720[1]), .C(n43564), .D(n19), 
         .Z(n790[1])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C+(D))+!B (C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_174_i2_4_lut.init = 16'h5c50;
    LUT4 i3614_3_lut_4_lut (.A(n429[2]), .B(n45807), .C(n429[1]), .D(n23471), 
         .Z(n6_adj_373)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !((C (D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3614_3_lut_4_lut.init = 16'h7331;
    LUT4 i38172_2_lut_rep_811_3_lut_4_lut_4_lut_4_lut_4_lut (.A(n45953), .B(n45946), 
         .C(n45975), .D(n45952), .Z(n45932)) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;
    defparam i38172_2_lut_rep_811_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h3323;
    LUT4 div_53_i155_3_lut_3_lut_3_lut_4_lut_4_lut_4_lut (.A(n45953), .B(n45938), 
         .C(n45954), .D(n45946), .Z(n222_adj_334)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;
    defparam div_53_i155_3_lut_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h4bf0;
    PFUMX i38368 (.BLUT(n45620), .ALUT(n45619), .C0(n45872), .Z(n43689));
    LUT4 oprand_3__bdd_4_lut_38270 (.A(n46875), .B(oprand[4]), .C(oprand[1]), 
         .D(oprand[2]), .Z(n114)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;
    defparam oprand_3__bdd_4_lut_38270.init = 16'h07c0;
    LUT4 div_53_i157_3_lut_rep_804_3_lut_4_lut_4_lut_4_lut_4_lut_4_lut (.A(n45953), 
         .B(n45946), .C(n45975), .D(n45952), .Z(n45925)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A (B (C (D)+!C !(D))+!B !(C+(D)))) */ ;
    defparam div_53_i157_3_lut_rep_804_3_lut_4_lut_4_lut_4_lut_4_lut_4_lut.init = 16'hc02f;
    CCU2D add_451_7 (.A0(n1842[4]), .B0(n1842[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40469), 
          .S0(n1855[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_451_7.INIT0 = 16'h5999;
    defparam add_451_7.INIT1 = 16'h0000;
    defparam add_451_7.INJECT1_0 = "NO";
    defparam add_451_7.INJECT1_1 = "NO";
    LUT4 i4774_4_lut (.A(n21777), .B(n45741), .C(n790[2]), .D(n45750), 
         .Z(n6_adj_485)) /* synthesis lut_function=(A+(B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i4774_4_lut.init = 16'heaae;
    LUT4 i15149_4_lut (.A(n9081), .B(n21776), .C(n43670), .D(n45757), 
         .Z(n21777)) /* synthesis lut_function=(!(A ((C (D)+!C !(D))+!B)+!A !(B (C (D)+!C !(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i15149_4_lut.init = 16'h4884;
    LUT4 i4773_4_lut (.A(n45741), .B(n790[1]), .C(n790[2]), .D(n45750), 
         .Z(n21776)) /* synthesis lut_function=(A+(B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i4773_4_lut.init = 16'heaae;
    LUT4 i1_2_lut_4_lut_adj_221 (.A(n43762), .B(n45833), .C(n43738), .D(n429[2]), 
         .Z(n4_adj_348)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_221.init = 16'h9669;
    LUT4 i2_4_lut_adj_222 (.A(n8_adj_486), .B(n45756), .C(n23070), .D(n4_adj_386), 
         .Z(n43673)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i2_4_lut_adj_222.init = 16'h6996;
    LUT4 i5246_4_lut (.A(n2476[3]), .B(n2476[5]), .C(n2476[2]), .D(n22479), 
         .Z(n8_adj_486)) /* synthesis lut_function=(A ((C (D))+!B)+!A !(B+!(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5246_4_lut.init = 16'hb232;
    LUT4 i2_4_lut_adj_223 (.A(n2476[5]), .B(n45752), .C(n45756), .D(n45740), 
         .Z(n7_adj_339)) /* synthesis lut_function=(!(A (B (C+(D)))+!A !(B (C+(D))))) */ ;
    defparam i2_4_lut_adj_223.init = 16'h666a;
    LUT4 i32142_2_lut_3_lut_4_lut (.A(n46183), .B(n9_adj_487), .C(oprand[0]), 
         .D(oprand[1]), .Z(n4)) /* synthesis lut_function=(A (B (C+!(D))+!B (C+(D)))+!A (C+!(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam i32142_2_lut_3_lut_4_lut.init = 16'hf2fd;
    CCU2D add_451_5 (.A0(n1842[2]), .B0(n1842[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1842[3]), .B1(n1842[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40468), .COUT(n40469), .S0(n1855[3]), .S1(n1855[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_451_5.INIT0 = 16'h5999;
    defparam add_451_5.INIT1 = 16'h5666;
    defparam add_451_5.INJECT1_0 = "NO";
    defparam add_451_5.INJECT1_1 = "NO";
    LUT4 mux_160_i2_3_lut (.A(n1855[5]), .B(n685[1]), .C(n89), .Z(n720[1])) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_160_i2_3_lut.init = 16'h5c5c;
    LUT4 i3_3_lut_4_lut (.A(n45808), .B(n41124), .C(n41282), .D(n43741), 
         .Z(n8_adj_372)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i3_3_lut_4_lut.init = 16'h9669;
    LUT4 div_53_i154_3_lut_3_lut_4_lut_4_lut_4_lut_4_lut (.A(n45961), .B(n191_adj_326), 
         .C(n45954), .D(n45945), .Z(n221_adj_333)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B (C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_i154_3_lut_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'hccc2;
    LUT4 i1_2_lut_3_lut_4_lut_adj_224 (.A(n46183), .B(n9_adj_487), .C(oprand[0]), 
         .D(oprand[1]), .Z(n41356)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam i1_2_lut_3_lut_4_lut_adj_224.init = 16'h2dd2;
    LUT4 i1_2_lut_rep_809_3_lut_4_lut (.A(n45985), .B(n45966), .C(n43353), 
         .D(n45944), .Z(n45930)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i1_2_lut_rep_809_3_lut_4_lut.init = 16'hf9f0;
    LUT4 i23898_2_lut_rep_657_3_lut_4_lut (.A(n46138), .B(n45783), .C(n46157), 
         .D(n45), .Z(n45778)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i23898_2_lut_rep_657_3_lut_4_lut.init = 16'h0080;
    LUT4 i32756_3_lut_4_lut (.A(n46188), .B(oprand[0]), .C(n46204), .D(n46170), 
         .Z(n12888[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam i32756_3_lut_4_lut.init = 16'h7f80;
    LUT4 i38101_4_lut (.A(n45780), .B(n45774), .C(n4_adj_488), .D(n45491), 
         .Z(n44729)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B (C (D))+!B (C+(D)))) */ ;
    defparam i38101_4_lut.init = 16'h84ed;
    CCU2D add_451_3 (.A0(n1842[0]), .B0(n1842[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1842[1]), .B1(n1842[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40467), .COUT(n40468), .S0(n1855[1]), .S1(n1855[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_451_3.INIT0 = 16'h5666;
    defparam add_451_3.INIT1 = 16'h5666;
    defparam add_451_3.INJECT1_0 = "NO";
    defparam add_451_3.INJECT1_1 = "NO";
    LUT4 div_39_i180_3_lut_rep_821_4_lut (.A(n45958), .B(n45957), .C(n18[2]), 
         .D(n45974), .Z(n45942)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_i180_3_lut_rep_821_4_lut.init = 16'hf1e0;
    LUT4 mux_174_i3_4_lut (.A(n2085[5]), .B(n45763), .C(n43564), .D(n19), 
         .Z(n790[2])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C+(D))+!B (C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_174_i3_4_lut.init = 16'h5c50;
    CCU2D add_451_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n45766), .B1(n40913), .C1(n46137), .D1(n650[1]), .COUT(n40467), 
          .S1(n1855[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_451_1.INIT0 = 16'hF000;
    defparam add_451_1.INIT1 = 16'h09f9;
    defparam add_451_1.INJECT1_0 = "NO";
    defparam add_451_1.INJECT1_1 = "NO";
    LUT4 mux_40_i3_3_lut_rep_823_4_lut (.A(n45958), .B(n45957), .C(n11), 
         .D(n45974), .Z(n45944)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_40_i3_3_lut_rep_823_4_lut.init = 16'hfe0e;
    LUT4 div_39_i174_3_lut_4_lut (.A(n45958), .B(n45957), .C(n18[8]), 
         .D(n45964), .Z(n250_adj_456)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_i174_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_146_i3_3_lut (.A(n1569[5]), .B(n615[2]), .C(n89_adj_303), 
         .Z(n650[2])) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_146_i3_3_lut.init = 16'h5c5c;
    LUT4 mux_139_i3_4_lut (.A(n43681), .B(n580[2]), .C(n46145), .D(n4_adj_489), 
         .Z(n615[2])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_139_i3_4_lut.init = 16'hc5ca;
    LUT4 div_39_i175_3_lut_4_lut (.A(n45958), .B(n45957), .C(n18[7]), 
         .D(n221), .Z(n251_adj_454)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_i175_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_225 (.A(n429[3]), .B(n45809), .C(n429[2]), 
         .D(n41124), .Z(n41354)) /* synthesis lut_function=(A (B (D)+!B (C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_3_lut_4_lut_adj_225.init = 16'hbd42;
    CCU2D add_449_7 (.A0(n1829[4]), .B0(n1829[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40466), 
          .S0(n1842[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_449_7.INIT0 = 16'h5999;
    defparam add_449_7.INIT1 = 16'h0000;
    defparam add_449_7.INJECT1_0 = "NO";
    defparam add_449_7.INJECT1_1 = "NO";
    LUT4 i5456_2_lut_rep_615_4_lut (.A(n2590[5]), .B(n895[4]), .C(n43563), 
         .D(n45749), .Z(n45736)) /* synthesis lut_function=(!(A (B (C (D))+!B (D))+!A !(B+(C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i5456_2_lut_rep_615_4_lut.init = 16'h5cff;
    LUT4 i3578_3_lut_4_lut (.A(n429[3]), .B(n45809), .C(n429[2]), .D(n41124), 
         .Z(n6_adj_466)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B ((D)+!C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3578_3_lut_4_lut.init = 16'h3173;
    CCU2D add_449_5 (.A0(n1829[2]), .B0(n1829[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1829[3]), .B1(n1829[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40465), .COUT(n40466), .S0(n1842[3]), .S1(n1842[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_449_5.INIT0 = 16'h5999;
    defparam add_449_5.INIT1 = 16'h5666;
    defparam add_449_5.INJECT1_0 = "NO";
    defparam add_449_5.INJECT1_1 = "NO";
    LUT4 i3923_4_lut (.A(n45795), .B(n45831), .C(n4_adj_396), .D(n45548), 
         .Z(n8_adj_490)) /* synthesis lut_function=(A (B (C (D))+!B (C+(D)))+!A !(B (C+!(D))+!B !((D)+!C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3923_4_lut.init = 16'hb721;
    LUT4 mux_132_i3_3_lut (.A(n1311[5]), .B(n545[2]), .C(n89_adj_320), 
         .Z(n580[2])) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_132_i3_3_lut.init = 16'h5c5c;
    CCU2D add_449_3 (.A0(n1829[0]), .B0(n1829[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1829[1]), .B1(n1829[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40464), .COUT(n40465), .S0(n1842[1]), .S1(n1842[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_449_3.INIT0 = 16'h5666;
    defparam add_449_3.INIT1 = 16'h5666;
    defparam add_449_3.INJECT1_0 = "NO";
    defparam add_449_3.INJECT1_1 = "NO";
    CCU2D add_449_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n6_adj_491), .B1(n5_adj_436), .C1(n46137), .D1(n650[2]), 
          .COUT(n40464), .S1(n1842[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_449_1.INIT0 = 16'hF000;
    defparam add_449_1.INIT1 = 16'h06f6;
    defparam add_449_1.INJECT1_0 = "NO";
    defparam add_449_1.INJECT1_1 = "NO";
    CCU2D add_447_7 (.A0(n1816[4]), .B0(n1816[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40463), 
          .S0(n1829[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_447_7.INIT0 = 16'h5999;
    defparam add_447_7.INIT1 = 16'h0000;
    defparam add_447_7.INJECT1_0 = "NO";
    defparam add_447_7.INJECT1_1 = "NO";
    LUT4 mux_146_i2_4_lut (.A(n1582[5]), .B(n580[1]), .C(n89_adj_303), 
         .D(n46145), .Z(n650[1])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C+(D))+!B (C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_146_i2_4_lut.init = 16'h5c50;
    LUT4 i1_2_lut_rep_688 (.A(n43714), .B(n43762), .Z(n45809)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_rep_688.init = 16'h6666;
    LUT4 i1_2_lut_rep_661 (.A(n23779), .B(n1687[5]), .Z(n45782)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_rep_661.init = 16'h6666;
    LUT4 mux_107_i4_3_lut_4_lut (.A(n43714), .B(n43762), .C(n37), .D(n429[3]), 
         .Z(n462[3])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_107_i4_3_lut_4_lut.init = 16'h6f60;
    LUT4 i3571_3_lut_rep_687_4_lut (.A(n43714), .B(n43762), .C(n429[2]), 
         .D(n429[3]), .Z(n45808)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C+!(D)))) */ ;
    defparam i3571_3_lut_rep_687_4_lut.init = 16'h90f9;
    LUT4 i2_3_lut_4_lut_adj_226 (.A(n43714), .B(n43762), .C(n429[3]), 
         .D(n429[2]), .Z(n23471)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i2_3_lut_4_lut_adj_226.init = 16'h6996;
    LUT4 i1_2_lut_4_lut_adj_227 (.A(n45994), .B(n45986), .C(n45960), .D(n45961), 
         .Z(n4_adj_325)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A (B (C+(D))+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_4_lut_adj_227.init = 16'hff6a;
    LUT4 i2_4_lut_adj_228 (.A(n45729), .B(n43706), .C(n45475), .D(n43647), 
         .Z(n6_adj_404)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;
    defparam i2_4_lut_adj_228.init = 16'h6c9c;
    LUT4 i5232_2_lut_4_lut (.A(n2358[5]), .B(n825[2]), .C(n45), .D(n45739), 
         .Z(n22479)) /* synthesis lut_function=(!(A (B (C (D))+!B (D))+!A !(B+(C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i5232_2_lut_4_lut.init = 16'h5cff;
    LUT4 mux_153_i4_3_lut_4_lut (.A(n23779), .B(n1687[5]), .C(n46137), 
         .D(n45790), .Z(n685[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam mux_153_i4_3_lut_4_lut.init = 16'hf909;
    LUT4 i5219_2_lut_4_lut (.A(n2358[5]), .B(n825[2]), .C(n45), .D(n2476[5]), 
         .Z(n2489[1])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(B (D)+!B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i5219_2_lut_4_lut.init = 16'ha35c;
    LUT4 i5856_2_lut_4_lut (.A(n43765), .B(n43732), .C(n45843), .D(n4_adj_380), 
         .Z(n21939)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C+(D)))) */ ;
    defparam i5856_2_lut_4_lut.init = 16'hff96;
    LUT4 i1_3_lut_4_lut_adj_229 (.A(n45743), .B(n45756), .C(n45738), .D(n2476[5]), 
         .Z(n23079)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_229.init = 16'h6966;
    LUT4 i1_2_lut_rep_620 (.A(n23806), .B(n43670), .Z(n45741)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_rep_620.init = 16'h6666;
    LUT4 mux_202_i2_4_lut (.A(n2629[5]), .B(n860[1]), .C(n43563), .D(n46157), 
         .Z(n930[1])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C+(D))+!B (C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_202_i2_4_lut.init = 16'h5c50;
    LUT4 i23996_4_lut (.A(n168), .B(n257), .C(n270_adj_514[1]), .D(n146[1]), 
         .Z(n30723)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C (D)))) */ ;
    defparam i23996_4_lut.init = 16'hfaee;
    LUT4 n43808_bdd_3_lut_4_lut_rep_835 (.A(n45973), .B(n45962), .C(n45966), 
         .D(n45972), .Z(n45956)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam n43808_bdd_3_lut_4_lut_rep_835.init = 16'h02fd;
    LUT4 mux_29_i1_4_lut (.A(n13_adj_492), .B(n159), .C(n7), .D(n45463), 
         .Z(n112[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_29_i1_4_lut.init = 16'hcfca;
    LUT4 i5_4_lut_adj_230 (.A(n159), .B(n10_adj_493), .C(n7_adj_494), 
         .D(n278_adj_495), .Z(n13_adj_492)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_230.init = 16'hfefc;
    LUT4 i2_3_lut_rep_645_4_lut (.A(n23779), .B(n1687[5]), .C(n40740), 
         .D(n44729), .Z(n45766)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i2_3_lut_rep_645_4_lut.init = 16'h6996;
    CCU2D add_447_5 (.A0(n1816[2]), .B0(n1816[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1816[3]), .B1(n1816[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40462), .COUT(n40463), .S0(n1829[3]), .S1(n1829[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_447_5.INIT0 = 16'h5999;
    defparam add_447_5.INIT1 = 16'h5666;
    defparam add_447_5.INJECT1_0 = "NO";
    defparam add_447_5.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_231 (.A(n15_adj_496), .B(n45980), .C(n261[2]), .D(n17[1]), 
         .Z(n10_adj_493)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_231.init = 16'hfaee;
    LUT4 i1_2_lut_4_lut_4_lut_adj_232 (.A(n45973), .B(n45962), .C(n45966), 
         .D(n45972), .Z(n6_adj_462)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B+(C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_4_lut_4_lut_adj_232.init = 16'h56ff;
    LUT4 i1_2_lut_rep_830_4_lut (.A(n45970), .B(n221), .C(n45964), .D(n45958), 
         .Z(n45951)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_rep_830_4_lut.init = 16'hfffe;
    CCU2D add_447_3 (.A0(n1816[0]), .B0(n1816[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1816[1]), .B1(n1816[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40461), .COUT(n40462), .S0(n1829[1]), .S1(n1829[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_447_3.INIT0 = 16'h5666;
    defparam add_447_3.INIT1 = 16'h5666;
    defparam add_447_3.INJECT1_0 = "NO";
    defparam add_447_3.INJECT1_1 = "NO";
    LUT4 div_39_i178_3_lut_4_lut_4_lut (.A(n45963), .B(n224), .C(n18[4]), 
         .D(n45957), .Z(n254_adj_453)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam div_39_i178_3_lut_4_lut_4_lut.init = 16'hf0c4;
    LUT4 div_28_i194_3_lut (.A(n246_adj_458), .B(n261[3]), .C(n17[1]), 
         .Z(n7_adj_494)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_i194_3_lut.init = 16'hcaca;
    LUT4 div_28_i196_3_lut (.A(n248), .B(n261[1]), .C(n17[1]), .Z(n278_adj_495)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_i196_3_lut.init = 16'hcaca;
    LUT4 i5855_2_lut_4_lut (.A(n43765), .B(n43732), .C(n45843), .D(n4_adj_380), 
         .Z(n9966)) /* synthesis lut_function=(A (B (C (D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C (D)))) */ ;
    defparam i5855_2_lut_4_lut.init = 16'h9600;
    CCU2D add_447_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n46870), .B1(n45782), .C1(n46144), .D1(n45790), .COUT(n40461), 
          .S1(n1829[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_447_1.INIT0 = 16'hF000;
    defparam add_447_1.INIT1 = 16'h04fe;
    defparam add_447_1.INJECT1_0 = "NO";
    defparam add_447_1.INJECT1_1 = "NO";
    CCU2D div_39_add_193_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n46264), .B1(n46266), .C1(n112[0]), .D1(n112[2]), 
          .COUT(n40410));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_add_193_1.INIT0 = 16'h0000;
    defparam div_39_add_193_1.INIT1 = 16'h0e1f;
    defparam div_39_add_193_1.INJECT1_0 = "NO";
    defparam div_39_add_193_1.INJECT1_1 = "NO";
    LUT4 div_28_i190_3_lut (.A(n242_adj_459), .B(n261[7]), .C(n17[1]), 
         .Z(n15_adj_496)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_i190_3_lut.init = 16'hcaca;
    LUT4 mux_181_i3_3_lut_4_lut (.A(n23806), .B(n43670), .C(n46138), .D(n790[2]), 
         .Z(n825[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam mux_181_i3_3_lut_4_lut.init = 16'hf909;
    LUT4 i1_4_lut_4_lut_adj_233 (.A(n23806), .B(n43670), .C(n6_adj_485), 
         .D(n40766), .Z(n43709)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C (D)))+!A !(B (C (D))+!B (C+(D))))) */ ;
    defparam i1_4_lut_4_lut_adj_233.init = 16'h533a;
    LUT4 mux_47_i3_3_lut_4_lut (.A(n45965), .B(n22712), .C(n46123), .D(n45944), 
         .Z(n73_adj_336)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A ((D)+!C)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_47_i3_3_lut_4_lut.init = 16'hfd0d;
    LUT4 div_46_i177_3_lut_rep_829_4_lut (.A(n45965), .B(n22712), .C(n45962), 
         .D(n45973), .Z(n45950)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (D))+!A (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_46_i177_3_lut_rep_829_4_lut.init = 16'h0df2;
    LUT4 i37208_4_lut (.A(n270_adj_514[6]), .B(n270_adj_514[7]), .C(n270_adj_514[5]), 
         .D(n270_adj_514[4]), .Z(n44099)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i37208_4_lut.init = 16'hfffe;
    LUT4 i37139_2_lut (.A(n270_adj_514[8]), .B(n270_adj_514[3]), .Z(n44026)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i37139_2_lut.init = 16'heeee;
    LUT4 i4479_3_lut_rep_654_4_lut (.A(n23779), .B(n1687[5]), .C(n6_adj_422), 
         .D(n40740), .Z(n45775)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C+!(D)))) */ ;
    defparam i4479_3_lut_rep_654_4_lut.init = 16'h90f9;
    LUT4 i37187_3_lut_rep_1050 (.A(n87), .B(n23565), .C(n4_adj_497), .Z(n46171)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i37187_3_lut_rep_1050.init = 16'hefef;
    LUT4 i37141_2_lut (.A(n18[8]), .B(n18[3]), .Z(n44028)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i37141_2_lut.init = 16'heeee;
    LUT4 i36957_2_lut (.A(n18[6]), .B(n18[5]), .Z(n43834)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i36957_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_234 (.A(n46225), .B(n109_adj_498), .C(akku_o_c_4), 
         .D(n8), .Z(n89_adj_320)) /* synthesis lut_function=(A (B ((D)+!C))+!A !((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_4_lut_adj_234.init = 16'h8c0c;
    LUT4 i1_4_lut_adj_235 (.A(n46345), .B(n46324), .C(n46330), .D(n46873), 
         .Z(n109_adj_498)) /* synthesis lut_function=(A (B (C))+!A !(((D)+!C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_4_lut_adj_235.init = 16'h80c0;
    CCU2D add_445_7 (.A0(n38301), .B0(n38297), .C0(n45878), .D0(n45879), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40460), 
          .S0(n1816[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_445_7.INIT0 = 16'h9a65;
    defparam add_445_7.INIT1 = 16'h0000;
    defparam add_445_7.INJECT1_0 = "NO";
    defparam add_445_7.INJECT1_1 = "NO";
    LUT4 i15757_2_lut_rep_668_4_lut (.A(n1829[5]), .B(n685[3]), .C(n89), 
         .D(n45791), .Z(n45789)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B (D)+!B ((D)+!C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i15757_2_lut_rep_668_4_lut.init = 16'h005c;
    CCU2D add_445_5 (.A0(n45818), .B0(n45892), .C0(n45822), .D0(n21753), 
          .A1(n45818), .B1(n4_adj_499), .C1(n21753), .D1(n23044), .CIN(n40459), 
          .COUT(n40460), .S0(n1816[3]), .S1(n1816[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_445_5.INIT0 = 16'ha659;
    defparam add_445_5.INIT1 = 16'h56a9;
    defparam add_445_5.INJECT1_0 = "NO";
    defparam add_445_5.INJECT1_1 = "NO";
    LUT4 i2_4_lut_rep_1162 (.A(n46019), .B(n46013), .C(n46081), .D(n6_adj_408), 
         .Z(n46848)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B (D)+!B !(D))) */ ;
    defparam i2_4_lut_rep_1162.init = 16'hc639;
    LUT4 i5443_2_lut_rep_614_4_lut_4_lut (.A(n43563), .B(n895[4]), .C(n2590[5]), 
         .Z(n45735)) /* synthesis lut_function=(A (C)+!A !(B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5443_2_lut_rep_614_4_lut_4_lut.init = 16'hb1b1;
    LUT4 i15039_3_lut_4_lut (.A(n45817), .B(n45815), .C(n41371), .D(n41285), 
         .Z(n21624)) /* synthesis lut_function=(!(A (D)+!A ((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i15039_3_lut_4_lut.init = 16'h00ae;
    CCU2D add_445_3 (.A0(n45879), .B0(n45820), .C0(n45822), .D0(GND_net), 
          .A1(n45879), .B1(n45820), .C1(n45822), .D1(n4400[0]), .CIN(n40458), 
          .COUT(n40459), .S0(n1816[1]), .S1(n1816[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_445_3.INIT0 = 16'h9969;
    defparam add_445_3.INIT1 = 16'h9669;
    defparam add_445_3.INJECT1_0 = "NO";
    defparam add_445_3.INJECT1_1 = "NO";
    CCU2D add_445_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n46870), .B1(n1687[5]), .C1(n46144), .D1(n45794), .COUT(n40458), 
          .S1(n1816[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_445_1.INIT0 = 16'hF000;
    defparam add_445_1.INIT1 = 16'h04fe;
    defparam add_445_1.INJECT1_0 = "NO";
    defparam add_445_1.INJECT1_1 = "NO";
    LUT4 i38135_2_lut_4_lut_4_lut (.A(n46240), .B(n4_adj_497), .C(n23565), 
         .D(n87), .Z(n43400)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i38135_2_lut_4_lut_4_lut.init = 16'hfff7;
    LUT4 i2_4_lut_adj_236 (.A(n46342), .B(oprand[0]), .C(n9_adj_487), 
         .D(n4_adj_500), .Z(n110)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i2_4_lut_adj_236.init = 16'hfefa;
    LUT4 mux_118_i6_4_lut (.A(n999[5]), .B(n462[5]), .C(n45_adj_356), 
         .D(n46196), .Z(n1156[2])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C+(D))+!B (C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_118_i6_4_lut.init = 16'h5c50;
    LUT4 mux_54_i5_3_lut_4_lut (.A(n160), .B(n45978), .C(n29_adj_353), 
         .D(n46001), .Z(n218[4])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam mux_54_i5_3_lut_4_lut.init = 16'hefe0;
    LUT4 n88_bdd_4_lut (.A(n46206), .B(akku_o_c_0), .C(n87_adj_314), .D(akku_o_c_1), 
         .Z(n45285)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)))+!A (B+(C+(D))))) */ ;
    defparam n88_bdd_4_lut.init = 16'h2801;
    LUT4 i1_2_lut_rep_1036_4_lut (.A(n46210), .B(n46209), .C(n46206), 
         .D(n43349), .Z(n46157)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_2_lut_rep_1036_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_1029_3_lut_3_lut (.A(n46271), .B(akku_o_c_1), .C(n46248), 
         .Z(n46150)) /* synthesis lut_function=(A (B+!(C))+!A (B (C)+!B !(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i1_2_lut_rep_1029_3_lut_3_lut.init = 16'hcbcb;
    CCU2D add_394_7 (.A0(n1569[4]), .B0(n1569[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40457), 
          .S0(n1582[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_394_7.INIT0 = 16'h5999;
    defparam add_394_7.INIT1 = 16'h0000;
    defparam add_394_7.INJECT1_0 = "NO";
    defparam add_394_7.INJECT1_1 = "NO";
    LUT4 i38131_2_lut_2_lut (.A(n31), .B(n43_adj_299), .Z(n11)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i38131_2_lut_2_lut.init = 16'h7777;
    LUT4 n4_bdd_4_lut (.A(n45911), .B(n4330[1]), .C(n22635), .D(n6_adj_419), 
         .Z(n866[4])) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;
    defparam n4_bdd_4_lut.init = 16'h1f78;
    LUT4 i54_4_lut_4_lut_3_lut (.A(n46271), .B(akku_o_c_1), .C(n46248), 
         .Z(n43)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;
    defparam i54_4_lut_4_lut_3_lut.init = 16'h8989;
    LUT4 i2_3_lut_rep_1058 (.A(n46876), .B(n23565), .C(akku_o_c_2), .Z(n46179)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(39[10:22])
    defparam i2_3_lut_rep_1058.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut_adj_237 (.A(oprand[2]), .B(n23565), .C(akku_o_c_2), 
         .D(n14), .Z(n5_adj_460)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(39[10:22])
    defparam i1_2_lut_4_lut_adj_237.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_adj_238 (.A(n46876), .B(n23565), .C(akku_o_c_2), 
         .D(n37_adj_318), .Z(n23650)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(39[10:22])
    defparam i1_2_lut_4_lut_adj_238.init = 16'h00fe;
    LUT4 akku_o_c_4_bdd_4_lut_38306_then_3_lut (.A(akku_o_c_1), .B(akku_o_c_2), 
         .C(akku_o_c_3), .Z(n46301)) /* synthesis lut_function=(!(A (B+(C))+!A (C))) */ ;
    defparam akku_o_c_4_bdd_4_lut_38306_then_3_lut.init = 16'h0707;
    LUT4 i2_4_lut_adj_239 (.A(n46844), .B(n46336), .C(n31179), .D(akku_o_c_4), 
         .Z(n45_adj_356)) /* synthesis lut_function=(!((B (C+(D))+!B (C))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i2_4_lut_adj_239.init = 16'h020a;
    LUT4 i2_3_lut_rep_825_4_lut (.A(n160), .B(n45978), .C(n45954), .D(n191_adj_326), 
         .Z(n45946)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i2_3_lut_rep_825_4_lut.init = 16'hfff8;
    LUT4 i1_3_lut_3_lut_rep_621_4_lut (.A(n2590[5]), .B(n895[4]), .C(n43563), 
         .D(n45749), .Z(n45742)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (D))+!A !(B (D)+!B (C (D)+!C !(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_3_lut_3_lut_rep_621_4_lut.init = 16'h5ca3;
    LUT4 i24451_4_lut (.A(n46195), .B(oprand[4]), .C(oprand[3]), .D(n6), 
         .Z(n31179)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam i24451_4_lut.init = 16'h444c;
    LUT4 i31606_2_lut_3_lut_4_lut (.A(n45971), .B(n45985), .C(n45972), 
         .D(n45973), .Z(n22[6])) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C)+!B !(C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i31606_2_lut_3_lut_4_lut.init = 16'hb40f;
    CCU2D add_394_5 (.A0(n1569[2]), .B0(n1569[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1569[3]), .B1(n1569[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40456), .COUT(n40457), .S0(n1582[3]), .S1(n1582[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_394_5.INIT0 = 16'h5999;
    defparam add_394_5.INIT1 = 16'h5666;
    defparam add_394_5.INJECT1_0 = "NO";
    defparam add_394_5.INJECT1_1 = "NO";
    LUT4 mux_202_i3_3_lut_rep_603 (.A(n2616[5]), .B(n895[2]), .C(n43563), 
         .Z(n45724)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_202_i3_3_lut_rep_603.init = 16'h5c5c;
    CCU2D add_1770_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40409), 
          .S0(akku_o_8__N_50[8]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(79[27:57])
    defparam add_1770_cout.INIT0 = 16'h0000;
    defparam add_1770_cout.INIT1 = 16'h0000;
    defparam add_1770_cout.INJECT1_0 = "NO";
    defparam add_1770_cout.INJECT1_1 = "NO";
    LUT4 n45691_bdd_4_lut (.A(n45691), .B(n46388), .C(n46873), .D(akku_o_c_4), 
         .Z(n45721)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n45691_bdd_4_lut.init = 16'hca00;
    LUT4 i15216_3_lut_4_lut (.A(n45729), .B(n45723), .C(n45725), .D(n23094), 
         .Z(n21872)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i15216_3_lut_4_lut.init = 16'h00fe;
    LUT4 i15020_3_lut_4_lut (.A(n41143), .B(n45816), .C(n41286), .D(n776[2]), 
         .Z(n21590)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i15020_3_lut_4_lut.init = 16'hef00;
    LUT4 i31619_2_lut_rep_820_3_lut_4_lut_4_lut (.A(n45972), .B(n221_adj_435), 
         .C(n45962), .D(n45973), .Z(n45941)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;
    defparam i31619_2_lut_rep_820_3_lut_4_lut_4_lut.init = 16'hfdff;
    CCU2D add_394_3 (.A0(n1569[0]), .B0(n1569[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1569[1]), .B1(n1569[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40455), .COUT(n40456), .S0(n1582[1]), .S1(n1582[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_394_3.INIT0 = 16'h5999;
    defparam add_394_3.INIT1 = 16'h5666;
    defparam add_394_3.INJECT1_0 = "NO";
    defparam add_394_3.INJECT1_1 = "NO";
    LUT4 i37105_2_lut_rep_662 (.A(n755[6]), .B(n43564), .Z(n45783)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i37105_2_lut_rep_662.init = 16'h2222;
    LUT4 akku_o_c_4_bdd_4_lut_38306_else_3_lut (.A(akku_o_c_1), .B(akku_o_c_2), 
         .C(akku_o_c_0), .D(akku_o_c_3), .Z(n46300)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;
    defparam akku_o_c_4_bdd_4_lut_38306_else_3_lut.init = 16'hec00;
    LUT4 div_46_i175_3_lut_4_lut_4_lut (.A(n45972), .B(n221_adj_435), .C(n45966), 
         .D(n45955), .Z(n251_adj_429)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B)) */ ;
    defparam div_46_i175_3_lut_4_lut_4_lut.init = 16'hccc6;
    LUT4 i5_4_lut_adj_240 (.A(n9_adj_478), .B(n117_adj_354), .C(n8_adj_394), 
         .D(n9), .Z(n43341)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i5_4_lut_adj_240.init = 16'hfffe;
    LUT4 i31611_2_lut_rep_828_3_lut_4_lut_4_lut (.A(n45972), .B(n45973), 
         .C(n45985), .D(n45971), .Z(n45949)) /* synthesis lut_function=(!(A (B ((D)+!C)))) */ ;
    defparam i31611_2_lut_rep_828_3_lut_4_lut_4_lut.init = 16'h77f7;
    LUT4 i5619_4_lut_4_lut (.A(n2371[2]), .B(n2371[5]), .C(n2371[1]), 
         .D(n2_adj_390), .Z(n6_adj_411)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5619_4_lut_4_lut.init = 16'heaa8;
    CCU2D add_394_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n46147), .B1(n9_adj_487), .C1(n43400), .D1(n580[1]), .COUT(n40455), 
          .S1(n1582[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_394_1.INIT0 = 16'hF000;
    defparam add_394_1.INIT1 = 16'h02ff;
    defparam add_394_1.INJECT1_0 = "NO";
    defparam add_394_1.INJECT1_1 = "NO";
    CCU2D add_392_7 (.A0(n1556[4]), .B0(n1556[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40454), 
          .S0(n1569[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_392_7.INIT0 = 16'h5999;
    defparam add_392_7.INIT1 = 16'h0000;
    defparam add_392_7.INJECT1_0 = "NO";
    defparam add_392_7.INJECT1_1 = "NO";
    LUT4 oprand_1__bdd_4_lut_38454 (.A(oprand[1]), .B(oprand[2]), .C(oprand[0]), 
         .D(n46193), .Z(n45404)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A (B (C+(D))+!B !(C (D))))) */ ;
    defparam oprand_1__bdd_4_lut_38454.init = 16'h1224;
    CCU2D add_392_5 (.A0(n1556[2]), .B0(n1556[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1556[3]), .B1(n1556[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40453), .COUT(n40454), .S0(n1569[3]), .S1(n1569[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_392_5.INIT0 = 16'h5999;
    defparam add_392_5.INIT1 = 16'h5666;
    defparam add_392_5.INJECT1_0 = "NO";
    defparam add_392_5.INJECT1_1 = "NO";
    LUT4 i38123_3_lut_rep_1006_4_lut_4_lut_4_lut (.A(n46156), .B(n46878), 
         .C(n78), .D(n43), .Z(n46127)) /* synthesis lut_function=(!(A (B (D))+!A !(B+(C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam i38123_3_lut_rep_1006_4_lut_4_lut_4_lut.init = 16'h76ff;
    CCU2D add_392_3 (.A0(n1556[0]), .B0(n1556[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1556[1]), .B1(n1556[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40452), .COUT(n40453), .S0(n1569[1]), .S1(n1569[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_392_3.INIT0 = 16'h5999;
    defparam add_392_3.INIT1 = 16'h5666;
    defparam add_392_3.INJECT1_0 = "NO";
    defparam add_392_3.INJECT1_1 = "NO";
    LUT4 i5498_2_lut_rep_605_3_lut_4_lut_4_lut_4_lut (.A(n46845), .B(n45749), 
         .C(n45728), .Z(n45726)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5498_2_lut_rep_605_3_lut_4_lut_4_lut_4_lut.init = 16'hf7f7;
    LUT4 pwr_bdd_2_lut_38322_rep_1024_3_lut_3_lut_4_lut (.A(akku_o_c_2), .B(n46213), 
         .C(n46212), .D(n45481), .Z(n46145)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;
    defparam pwr_bdd_2_lut_38322_rep_1024_3_lut_3_lut_4_lut.init = 16'hfff6;
    LUT4 i1_3_lut_rep_1039_4_lut (.A(akku_o_c_2), .B(n46213), .C(akku_o_c_1), 
         .D(n87), .Z(n46160)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_3_lut_rep_1039_4_lut.init = 16'hf600;
    LUT4 i1_3_lut_rep_1062 (.A(n4_adj_497), .B(n46212), .C(oprand[1]), 
         .Z(n46183)) /* synthesis lut_function=(A+!(B+(C))) */ ;
    defparam i1_3_lut_rep_1062.init = 16'habab;
    LUT4 i23890_2_lut_rep_1038_4_lut (.A(n4_adj_497), .B(n46212), .C(oprand[1]), 
         .D(n9_adj_487), .Z(n46159)) /* synthesis lut_function=(!(A (D)+!A (B+(C+(D))))) */ ;
    defparam i23890_2_lut_rep_1038_4_lut.init = 16'h00ab;
    LUT4 i57_3_lut_4_lut_3_lut (.A(n4_adj_497), .B(n46878), .C(n9_adj_487), 
         .Z(n31_adj_501)) /* synthesis lut_function=(!(A (B+(C))+!A !(B))) */ ;
    defparam i57_3_lut_4_lut_3_lut.init = 16'h4646;
    LUT4 rem_66_i98_3_lut_4_lut_4_lut (.A(n4_adj_497), .B(n46212), .C(oprand[1]), 
         .D(n9_adj_487), .Z(n106)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+!(D)))+!A (B (C)+!B !(C+!(D)))) */ ;
    defparam rem_66_i98_3_lut_4_lut_4_lut.init = 16'hc3c8;
    LUT4 i3547_2_lut_4_lut_3_lut_4_lut (.A(n45817), .B(n429[3]), .C(n45841), 
         .D(n41371), .Z(n7658)) /* synthesis lut_function=(A (B+!(C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3547_2_lut_4_lut_3_lut_4_lut.init = 16'h8aaa;
    LUT4 i38435_then_4_lut (.A(oprand[1]), .B(oprand[0]), .C(oprand[3]), 
         .D(oprand[4]), .Z(n46864)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i38435_then_4_lut.init = 16'h0040;
    LUT4 i37241_2_lut_3_lut_4_lut (.A(n755[6]), .B(n43564), .C(n45), .D(n46138), 
         .Z(n30)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i37241_2_lut_3_lut_4_lut.init = 16'hfdff;
    LUT4 i1_3_lut_4_lut_4_lut_adj_241 (.A(n45745), .B(n45736), .C(n45747), 
         .Z(n7_adj_406)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_3_lut_4_lut_4_lut_adj_241.init = 16'h5656;
    LUT4 i1_2_lut_adj_242 (.A(n39_adj_313), .B(n51_adj_345), .Z(n37)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_2_lut_adj_242.init = 16'h8888;
    LUT4 rem_50_i76_3_lut_3_lut_4_lut (.A(n46206), .B(akku_o_c_1), .C(n86), 
         .D(n87_adj_314), .Z(n7_adj_502)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam rem_50_i76_3_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 i1_2_lut_rep_618_4_lut (.A(n2345[5]), .B(n825[3]), .C(n45), .D(n45756), 
         .Z(n45739)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(B (D)+!B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_618_4_lut.init = 16'ha35c;
    LUT4 i33683_2_lut_4_lut_4_lut (.A(n46206), .B(akku_o_c_1), .C(n86), 
         .D(n87_adj_314), .Z(n107_adj_503)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C))+!A (B (C)+!B !(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i33683_2_lut_4_lut_4_lut.init = 16'h343c;
    LUT4 rem_50_i77_3_lut_4_lut (.A(n46206), .B(akku_o_c_1), .C(n86), 
         .D(n87_adj_314), .Z(n106_adj_504)) /* synthesis lut_function=(!(A (B (C+(D)))+!A !(B (C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam rem_50_i77_3_lut_4_lut.init = 16'h626a;
    LUT4 i3542_4_lut_rep_691_4_lut (.A(n45817), .B(n429[3]), .C(n45841), 
         .D(n41371), .Z(n45812)) /* synthesis lut_function=(A (B+!(C (D)))+!A !((C+(D))+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3542_4_lut_rep_691_4_lut.init = 16'h8aae;
    LUT4 i37114_2_lut_rep_658_3_lut_4_lut (.A(n755[6]), .B(n43564), .C(n45), 
         .D(n46138), .Z(n45779)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i37114_2_lut_rep_658_3_lut_4_lut.init = 16'h0200;
    LUT4 i5_3_lut_4_lut (.A(n46270), .B(akku_o_c_1), .C(n46870), .D(n9_adj_484), 
         .Z(n14_adj_439)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i5_3_lut_4_lut.init = 16'hfff4;
    LUT4 i8_4_lut (.A(n15_adj_505), .B(n30175), .C(n14_adj_506), .D(n30180), 
         .Z(n15_adj_316)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i8_4_lut.init = 16'hfffe;
    LUT4 i14906_3_lut_4_lut (.A(n46054), .B(n46027), .C(n45979), .D(n23445), 
         .Z(n21411)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i14906_3_lut_4_lut.init = 16'h00fd;
    LUT4 i2_3_lut_4_lut_adj_243 (.A(n45817), .B(n429[3]), .C(n45841), 
         .D(n41371), .Z(n41282)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_4_lut_adj_243.init = 16'h24db;
    LUT4 i5197_2_lut_rep_619_4_lut (.A(n2345[5]), .B(n825[3]), .C(n45), 
         .D(n45758), .Z(n45740)) /* synthesis lut_function=(!(A (B (C (D))+!B (D))+!A !(B+(C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i5197_2_lut_rep_619_4_lut.init = 16'h5cff;
    LUT4 i6_4_lut_adj_244 (.A(n106_adj_504), .B(n107_adj_503), .C(n114), 
         .D(n46186), .Z(n15_adj_505)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i6_4_lut_adj_244.init = 16'hfffe;
    LUT4 div_39_i153_3_lut_rep_843_4_lut (.A(n191), .B(n45983), .C(n45992), 
         .D(n190), .Z(n45964)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_i153_3_lut_rep_843_4_lut.init = 16'hfe01;
    LUT4 i1_2_lut_4_lut_adj_245 (.A(n45817), .B(n429[3]), .C(n45841), 
         .D(n41285), .Z(n6_adj_470)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_4_lut_adj_245.init = 16'h718e;
    LUT4 i5_4_lut_adj_246 (.A(n7_adj_502), .B(n30168), .C(n46318), .D(n46870), 
         .Z(n14_adj_506)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i5_4_lut_adj_246.init = 16'hfffe;
    LUT4 i2_3_lut_4_lut_adj_247 (.A(n45819), .B(n45842), .C(n363[2]), 
         .D(n41388), .Z(n22740)) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_4_lut_adj_247.init = 16'hdb24;
    LUT4 i3_3_lut_rep_836_4_lut (.A(n45989), .B(n45981), .C(n45964), .D(n221), 
         .Z(n45957)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_3_lut_rep_836_4_lut.init = 16'hfffe;
    LUT4 i3157_3_lut_4_lut (.A(n45819), .B(n45842), .C(n363[2]), .D(n41388), 
         .Z(n6_adj_378)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (B (C (D))+!B (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3157_3_lut_4_lut.init = 16'h04df;
    LUT4 i24058_2_lut_4_lut (.A(n45819), .B(n363[2]), .C(n37_adj_301), 
         .D(n41286), .Z(n30785)) /* synthesis lut_function=(A (B+(C+!(D)))+!A !(B (C (D))+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i24058_2_lut_4_lut.init = 16'hacff;
    LUT4 i3299_2_lut_rep_693_4_lut (.A(n45819), .B(n363[2]), .C(n37_adj_301), 
         .D(n41143), .Z(n45814)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B ((D)+!C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i3299_2_lut_rep_693_4_lut.init = 16'hffac;
    LUT4 i1_2_lut_rep_696 (.A(n866[4]), .B(n43714), .Z(n45817)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_rep_696.init = 16'h6666;
    LUT4 i3535_4_lut_rep_694_4_lut (.A(n866[4]), .B(n43714), .C(n45841), 
         .D(n429[3]), .Z(n45815)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C+!(D))))) */ ;
    defparam i3535_4_lut_rep_694_4_lut.init = 16'h6f06;
    LUT4 i23762_2_lut_rep_844_3_lut (.A(n46009), .B(n46849), .C(n45985), 
         .Z(n45965)) /* synthesis lut_function=(!(A (B (C))+!A !(B+!(C)))) */ ;
    defparam i23762_2_lut_rep_844_3_lut.init = 16'h6f6f;
    LUT4 i2_3_lut_rep_930_4_lut (.A(n46067), .B(n37), .C(n22585), .D(n46136), 
         .Z(n46051)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i2_3_lut_rep_930_4_lut.init = 16'h2000;
    LUT4 mux_107_i5_3_lut_4_lut (.A(n866[4]), .B(n43714), .C(n37), .D(n45841), 
         .Z(n462[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;
    defparam mux_107_i5_3_lut_4_lut.init = 16'h9f90;
    CCU2D add_1770_9 (.A0(GND_net), .B0(n46133), .C0(n45771), .D0(akku_o_c_6), 
          .A1(GND_net), .B1(n46133), .C1(n46018), .D1(akku_o_c_7), .CIN(n40408), 
          .COUT(n40409), .S0(akku_o_8__N_50[6]), .S1(akku_o_8__N_50[7]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(79[27:57])
    defparam add_1770_9.INIT0 = 16'h596a;
    defparam add_1770_9.INIT1 = 16'h596a;
    defparam add_1770_9.INJECT1_0 = "NO";
    defparam add_1770_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_761_4_lut_4_lut (.A(n46019), .B(n46013), .C(n46081), 
         .D(n6_adj_408), .Z(n45882)) /* synthesis lut_function=(A (B (D)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;
    defparam i1_2_lut_rep_761_4_lut_4_lut.init = 16'hf807;
    LUT4 i1_2_lut_rep_827_3_lut_3_lut_4_lut (.A(n46009), .B(n46849), .C(n22712), 
         .D(n45985), .Z(n45948)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;
    defparam i1_2_lut_rep_827_3_lut_3_lut_4_lut.init = 16'hf90f;
    LUT4 i31593_2_lut_rep_841_3_lut (.A(n46009), .B(n46849), .C(n45985), 
         .Z(n45962)) /* synthesis lut_function=(A (B (C))+!A !(B+!(C))) */ ;
    defparam i31593_2_lut_rep_841_3_lut.init = 16'h9090;
    LUT4 i38435_else_4_lut (.A(oprand[1]), .B(oprand[0]), .C(oprand[3]), 
         .D(oprand[4]), .Z(n46863)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+(C+(D))))) */ ;
    defparam i38435_else_4_lut.init = 16'h2001;
    PFUMX i38357 (.BLUT(n45596), .ALUT(n396[7]), .C0(n45917), .Z(n43750));
    LUT4 i24103_2_lut_rep_845_4_lut (.A(n46009), .B(n46849), .C(n22712), 
         .D(n45985), .Z(n45966)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C))+!A (B (C)+!B (C+(D))))) */ ;
    defparam i24103_2_lut_rep_845_4_lut.init = 16'h060f;
    LUT4 mux_111_i2_3_lut_4_lut (.A(n46230), .B(n46229), .C(n462[1]), 
         .D(n45859), .Z(n475[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(39[10:22])
    defparam mux_111_i2_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i38348 (.BLUT(n45571), .ALUT(n45570), .C0(n583), .Z(n45572));
    LUT4 i1_3_lut_adj_248 (.A(akku_o_c_3), .B(akku_o_c_2), .C(akku_o_c_4), 
         .Z(n87_adj_314)) /* synthesis lut_function=(!((B (C))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i1_3_lut_adj_248.init = 16'h2a2a;
    CCU2D add_392_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n43681), .B1(n4_adj_489), .C1(n46145), .D1(n580[2]), .COUT(n40452), 
          .S1(n1569[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_392_1.INIT0 = 16'hF000;
    defparam add_392_1.INIT1 = 16'h09f9;
    defparam add_392_1.INJECT1_0 = "NO";
    defparam add_392_1.INJECT1_1 = "NO";
    LUT4 i37225_2_lut_rep_775_3_lut_4_lut (.A(n46230), .B(n46229), .C(n45_adj_356), 
         .D(n45904), .Z(n45896)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(39[10:22])
    defparam i37225_2_lut_rep_775_3_lut_4_lut.init = 16'h0e00;
    LUT4 mux_111_i1_3_lut_4_lut (.A(n46230), .B(n46229), .C(n462[0]), 
         .D(n462[4]), .Z(n475[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(39[10:22])
    defparam mux_111_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2_3_lut_4_lut_adj_249 (.A(n866[4]), .B(n43714), .C(n45841), 
         .D(n429[3]), .Z(n41124)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i2_3_lut_4_lut_adj_249.init = 16'h6996;
    LUT4 n1701_bdd_3_lut_4_lut_4_lut (.A(n45790), .B(n1687[5]), .C(n650[2]), 
         .D(n23779), .Z(n45490)) /* synthesis lut_function=(A (B (C (D))+!B !(C+!(D)))+!A !(B (C+(D))+!B ((D)+!C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam n1701_bdd_3_lut_4_lut_4_lut.init = 16'h8214;
    LUT4 div_46_i178_4_lut_3_lut_3_lut_4_lut (.A(n46009), .B(n46849), .C(n22712), 
         .D(n45985), .Z(n254_adj_430)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B (C (D))+!B !(D)))) */ ;
    defparam div_46_i178_4_lut_3_lut_3_lut_4_lut.init = 16'h6099;
    LUT4 i2013_3_lut_4_lut (.A(address[3]), .B(n46237), .C(address[4]), 
         .D(address[5]), .Z(pc_5__N_35[5])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i2013_3_lut_4_lut.init = 16'h7f80;
    LUT4 i4699_2_lut_rep_638_3_lut_4_lut_4_lut_3_lut (.A(n45789), .B(n45787), 
         .C(n45761), .Z(n45759)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i4699_2_lut_rep_638_3_lut_4_lut_4_lut_3_lut.init = 16'he0e0;
    LUT4 mux_160_i6_3_lut_4_lut (.A(n45879), .B(n45820), .C(n89), .D(n45822), 
         .Z(n720[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_160_i6_3_lut_4_lut.init = 16'h9f90;
    CCU2D add_1770_7 (.A0(address[4]), .B0(n46133), .C0(n46845), .D0(akku_o_c_4), 
          .A1(GND_net), .B1(n46133), .C1(n45749), .D1(akku_o_c_5), .CIN(n40407), 
          .COUT(n40408), .S0(akku_o_8__N_50[4]), .S1(akku_o_8__N_50[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(79[27:57])
    defparam add_1770_7.INIT0 = 16'hd1e2;
    defparam add_1770_7.INIT1 = 16'h596a;
    defparam add_1770_7.INJECT1_0 = "NO";
    defparam add_1770_7.INJECT1_1 = "NO";
    LUT4 i31603_2_lut_rep_834_3_lut_4_lut_4_lut (.A(n46000), .B(n46009), 
         .C(n46849), .D(n45985), .Z(n45955)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+!(D)))+!A ((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i31603_2_lut_rep_834_3_lut_4_lut_4_lut.init = 16'hdb59;
    LUT4 i1_3_lut_4_lut_adj_250 (.A(n46875), .B(n46233), .C(oprand[4]), 
         .D(n46305), .Z(n103)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam i1_3_lut_4_lut_adj_250.init = 16'hef00;
    LUT4 i23989_2_lut_rep_842_4_lut (.A(n112[4]), .B(n112[2]), .C(n46207), 
         .D(n45982), .Z(n45963)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i23989_2_lut_rep_842_4_lut.init = 16'hcaff;
    LUT4 i32749_2_lut_3_lut_4_lut_4_lut (.A(oprand[2]), .B(n46257), .C(oprand[1]), 
         .D(oprand[0]), .Z(n12888[2])) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A !(B (C)+!B (C (D))))) */ ;
    defparam i32749_2_lut_3_lut_4_lut_4_lut.init = 16'h5a6a;
    PFUMX i38346 (.BLUT(n45568), .ALUT(n45567), .C0(n41077), .Z(n41385));
    LUT4 i2_3_lut_rep_1056_4_lut (.A(akku_o_c_2), .B(n46258), .C(n46209), 
         .D(n46210), .Z(n46177)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (C+(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i2_3_lut_rep_1056_4_lut.init = 16'hfff2;
    LUT4 n88_bdd_3_lut_4_lut (.A(akku_o_c_2), .B(n46258), .C(akku_o_c_1), 
         .D(akku_o_c_0), .Z(n45284)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam n88_bdd_3_lut_4_lut.init = 16'h0200;
    LUT4 mux_33_i4_3_lut_rep_887_4_lut (.A(n46266), .B(n46264), .C(n112[3]), 
         .D(n112[5]), .Z(n46008)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam mux_33_i4_3_lut_rep_887_4_lut.init = 16'hf1e0;
    LUT4 i7821_1_lut_3_lut_4_lut (.A(n46266), .B(n46264), .C(n112[3]), 
         .D(n112[5]), .Z(n8_adj_451)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i7821_1_lut_3_lut_4_lut.init = 16'h0e1f;
    LUT4 mux_33_i5_3_lut_rep_929_4_lut (.A(n46266), .B(n46264), .C(n112[4]), 
         .D(n112[6]), .Z(n46050)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam mux_33_i5_3_lut_rep_929_4_lut.init = 16'hf1e0;
    LUT4 mux_33_i3_3_lut_rep_853_4_lut (.A(n46266), .B(n46264), .C(n112[2]), 
         .D(n112[4]), .Z(n45974)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam mux_33_i3_3_lut_rep_853_4_lut.init = 16'hf1e0;
    CCU2D add_390_7 (.A0(n1543[4]), .B0(n1543[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40451), 
          .S0(n1556[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_390_7.INIT0 = 16'h5999;
    defparam add_390_7.INIT1 = 16'h0000;
    defparam add_390_7.INJECT1_0 = "NO";
    defparam add_390_7.INJECT1_1 = "NO";
    LUT4 mux_33_i2_3_lut_4_lut (.A(n46266), .B(n46264), .C(n112[1]), .D(n112[3]), 
         .Z(n257)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam mux_33_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_33_i1_3_lut_4_lut (.A(n46266), .B(n46264), .C(n112[0]), .D(n112[2]), 
         .Z(n168)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam mux_33_i1_3_lut_4_lut.init = 16'hf1e0;
    CCU2D add_390_5 (.A0(n1543[2]), .B0(n1543[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1543[3]), .B1(n1543[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40450), .COUT(n40451), .S0(n1556[3]), .S1(n1556[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_390_5.INIT0 = 16'h5999;
    defparam add_390_5.INIT1 = 16'h5666;
    defparam add_390_5.INJECT1_0 = "NO";
    defparam add_390_5.INJECT1_1 = "NO";
    LUT4 div_53_i133_3_lut_4_lut_3_lut_4_lut (.A(n45994), .B(n45986), .C(n160), 
         .D(n161_adj_302), .Z(n191_adj_326)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A !((D)+!C)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_i133_3_lut_4_lut_3_lut_4_lut.init = 16'h8870;
    CCU2D add_390_3 (.A0(n1543[0]), .B0(n1543[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1543[1]), .B1(n1543[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40449), .COUT(n40450), .S0(n1556[1]), .S1(n1556[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_390_3.INIT0 = 16'h5999;
    defparam add_390_3.INIT1 = 16'h5666;
    defparam add_390_3.INJECT1_0 = "NO";
    defparam add_390_3.INJECT1_1 = "NO";
    LUT4 i132_then_4_lut_adj_251 (.A(akku_o_c_3), .B(akku_o_c_1), .C(akku_o_c_4), 
         .D(akku_o_c_2), .Z(n46304)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i132_then_4_lut_adj_251.init = 16'h1000;
    LUT4 i1_2_lut_4_lut_adj_252 (.A(n43732), .B(n41291), .C(n45850), .D(n363[2]), 
         .Z(n4_adj_379)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_252.init = 16'h9669;
    CCU2D add_390_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n6_adj_399), .B1(n5_adj_507), .C1(n46145), .D1(n45799), 
          .COUT(n40449), .S1(n1556[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_390_1.INIT0 = 16'hF000;
    defparam add_390_1.INIT1 = 16'h06f6;
    defparam add_390_1.INJECT1_0 = "NO";
    defparam add_390_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_253 (.A(oprand[2]), .B(n46245), .C(n46258), 
         .D(akku_o_c_2), .Z(n8_adj_338)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam i1_2_lut_3_lut_4_lut_adj_253.init = 16'h8f88;
    LUT4 i20_4_lut_4_lut_3_lut (.A(\states[1] ), .B(states[0]), .C(states_c[2]), 
         .Z(clk_c_enable_20)) /* synthesis lut_function=(!(A (B)+!A !(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam i20_4_lut_4_lut_3_lut.init = 16'h7272;
    LUT4 i2_2_lut_rep_839_3_lut_4_lut (.A(n45994), .B(n45986), .C(n160), 
         .D(n161_adj_302), .Z(n45960)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_2_lut_rep_839_3_lut_4_lut.init = 16'hfff8;
    LUT4 i36987_3_lut_2_lut_rep_840_3_lut_4_lut (.A(n45994), .B(n45986), 
         .C(n160), .D(n161_adj_302), .Z(n45961)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i36987_3_lut_2_lut_rep_840_3_lut_4_lut.init = 16'hf080;
    LUT4 i15124_3_lut_rep_659_4_lut_4_lut (.A(n45790), .B(n1687[5]), .C(n650[2]), 
         .D(n23779), .Z(n45780)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A !(B (C+(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i15124_3_lut_rep_659_4_lut_4_lut.init = 16'h6462;
    LUT4 i2_3_lut_rep_664 (.A(n1687[5]), .B(n45794), .C(n45790), .Z(n45785)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;
    defparam i2_3_lut_rep_664.init = 16'hc6c6;
    LUT4 i1_2_lut_3_lut_4_lut_adj_254 (.A(n1687[5]), .B(n45794), .C(n45790), 
         .D(n23779), .Z(n4_adj_488)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B !(D))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_254.init = 16'h936c;
    LUT4 div_53_i134_3_lut_rep_833_4_lut_4_lut (.A(n45994), .B(n45986), 
         .C(n161_adj_302), .D(n160), .Z(n45954)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_53_i134_3_lut_rep_833_4_lut_4_lut.init = 16'h6662;
    LUT4 i1_2_lut_adj_255 (.A(n39_adj_343), .B(n51_adj_344), .Z(n37_adj_301)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_2_lut_adj_255.init = 16'h8888;
    LUT4 i24149_2_lut_4_lut (.A(n217), .B(n231[2]), .C(n45991), .D(n248), 
         .Z(n30876)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i24149_2_lut_4_lut.init = 16'hca00;
    LUT4 i23992_2_lut_rep_837_3_lut_4_lut (.A(n46008), .B(n45992), .C(n224), 
         .D(n45974), .Z(n45958)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (B (C (D))+!B (C))) */ ;
    defparam i23992_2_lut_rep_837_3_lut_4_lut.init = 16'hf090;
    LUT4 i4_4_lut_adj_256 (.A(n7_adj_322), .B(n46156), .C(n23565), .D(n78), 
         .Z(n15)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i4_4_lut_adj_256.init = 16'hfffe;
    LUT4 i37143_2_lut_4_lut_4_lut (.A(n46008), .B(n45992), .C(n45969), 
         .D(n190), .Z(n44030)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A ((D)+!B)) */ ;
    defparam i37143_2_lut_4_lut_4_lut.init = 16'hfd9b;
    LUT4 i1_3_lut_4_lut_adj_257 (.A(n46268), .B(akku_o_c_4), .C(n46367), 
         .D(n46859), .Z(n110_adj_311)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_257.init = 16'hfff4;
    LUT4 i1_3_lut_4_lut_adj_258 (.A(oprand[4]), .B(n46250), .C(n45374), 
         .D(n46264), .Z(n43554)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_3_lut_4_lut_adj_258.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_259 (.A(n46790), .B(n46876), .C(n46167), 
         .D(n46869), .Z(n37_adj_318)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_259.init = 16'h0200;
    LUT4 i2_2_lut_3_lut_4_lut_4_lut (.A(n45889), .B(n45823), .C(n23779), 
         .D(n45794), .Z(n6_adj_491)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(B (C)+!B (C (D)+!C !(D)))) */ ;
    defparam i2_2_lut_3_lut_4_lut_4_lut.init = 16'ha596;
    LUT4 div_39_i154_3_lut_4_lut (.A(n46005), .B(n45988), .C(n45992), 
         .D(n191), .Z(n221)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_i154_3_lut_4_lut.init = 16'hfe01;
    LUT4 i15118_2_lut_rep_672_4_lut_4_lut (.A(n45829), .B(n89_adj_303), 
         .C(n615[4]), .D(n1543[5]), .Z(n45793)) /* synthesis lut_function=(!(A ((D)+!B)+!A (B (D)+!B !(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i15118_2_lut_rep_672_4_lut_4_lut.init = 16'h10dc;
    LUT4 i4_2_lut_3_lut_4_lut (.A(oprand[4]), .B(n46256), .C(n117_adj_323), 
         .D(oprand[1]), .Z(n13)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C+(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam i4_2_lut_3_lut_4_lut.init = 16'hf7f0;
    LUT4 i32742_2_lut_3_lut_4_lut (.A(oprand[4]), .B(n46256), .C(oprand[0]), 
         .D(oprand[1]), .Z(n12888[1])) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam i32742_2_lut_3_lut_4_lut.init = 16'h87f0;
    LUT4 i2_4_lut_else_4_lut_adj_260 (.A(akku_o_c_0), .B(akku_o_c_4), .C(akku_o_c_2), 
         .D(akku_o_c_3), .Z(n46857)) /* synthesis lut_function=(!((B (C+!(D))+!B ((D)+!C))+!A)) */ ;
    defparam i2_4_lut_else_4_lut_adj_260.init = 16'h0820;
    CCU2D add_388_7 (.A0(VCC_net), .B0(n6_adj_369), .C0(n46045), .D0(n4_adj_403), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40448), 
          .S0(n1543[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_388_7.INIT0 = 16'ha995;
    defparam add_388_7.INIT1 = 16'h0000;
    defparam add_388_7.INJECT1_0 = "NO";
    defparam add_388_7.INJECT1_1 = "NO";
    LUT4 i1_4_lut_rep_1163 (.A(n45997), .B(n191_adj_335), .C(n12_adj_508), 
         .Z(n46849)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_4_lut_rep_1163.init = 16'h1010;
    LUT4 mux_202_i4_3_lut_rep_607 (.A(n2603[5]), .B(n895[3]), .C(n43563), 
         .Z(n45728)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_202_i4_3_lut_rep_607.init = 16'h5c5c;
    LUT4 i1_2_lut_rep_671_3_lut_3_lut_4_lut (.A(n45829), .B(n89_adj_303), 
         .C(n45794), .D(n45889), .Z(n45792)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (D))+!A (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_671_3_lut_3_lut_4_lut.init = 16'h0df2;
    LUT4 i31666_2_lut_rep_848_3_lut_4_lut (.A(n46007), .B(n45996), .C(n191), 
         .D(n46005), .Z(n45969)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i31666_2_lut_rep_848_3_lut_4_lut.init = 16'hfff8;
    CCU2D add_388_5 (.A0(VCC_net), .B0(n45829), .C0(n23019), .D0(n45887), 
          .A1(n1530[3]), .B1(n6_adj_369), .C1(n4_adj_403), .D1(n46045), 
          .CIN(n40447), .COUT(n40448), .S0(n1543[3]), .S1(n1543[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_388_5.INIT0 = 16'ha569;
    defparam add_388_5.INIT1 = 16'h5555;
    defparam add_388_5.INJECT1_0 = "NO";
    defparam add_388_5.INJECT1_1 = "NO";
    CCU2D add_388_3 (.A0(n45829), .B0(n4233[3]), .C0(n38213), .D0(n22463), 
          .A1(n40970), .B1(n6_adj_369), .C1(n4_adj_403), .D1(n46045), 
          .CIN(n40446), .COUT(n40447), .S0(n1543[1]), .S1(n1543[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_388_3.INIT0 = 16'ha956;
    defparam add_388_3.INIT1 = 16'h5555;
    defparam add_388_3.INJECT1_0 = "NO";
    defparam add_388_3.INJECT1_1 = "NO";
    LUT4 div_39_i155_3_lut_4_lut_rep_868 (.A(n46007), .B(n45996), .C(n45992), 
         .D(n46005), .Z(n45989)) /* synthesis lut_function=(A (B (D)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_i155_3_lut_4_lut_rep_868.init = 16'hf807;
    LUT4 i36950_2_lut_rep_849_4_lut_4_lut (.A(n46007), .B(n45996), .C(n45992), 
         .D(n46005), .Z(n45970)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i36950_2_lut_rep_849_4_lut_4_lut.init = 16'hfea7;
    LUT4 i31550_2_lut_3_lut_4_lut (.A(n45829), .B(n89_adj_303), .C(n45892), 
         .D(n46137), .Z(n4_adj_499)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i31550_2_lut_3_lut_4_lut.init = 16'h2f0f;
    PFUMX i38762 (.BLUT(n46863), .ALUT(n46864), .C0(n46876), .Z(n39_adj_343));
    LUT4 i1_2_lut_3_lut_4_lut_adj_261 (.A(n45829), .B(n89_adj_303), .C(n45885), 
         .D(n45889), .Z(n22896)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A (C)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_3_lut_4_lut_adj_261.init = 16'hf0d2;
    LUT4 div_28_i169_3_lut_4_lut (.A(n46004), .B(n22716), .C(n231[7]), 
         .D(n212), .Z(n242_adj_459)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_i169_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_28_i168_3_lut_4_lut (.A(n46004), .B(n22716), .C(n231[8]), 
         .D(n211), .Z(n241)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_i168_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_28_i170_3_lut_4_lut (.A(n46004), .B(n22716), .C(n231[6]), 
         .D(n213), .Z(n243)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_i170_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_28_i172_3_lut_4_lut (.A(n46004), .B(n22716), .C(n231[4]), 
         .D(n215), .Z(n245)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_i172_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15777_2_lut_3_lut_4_lut_4_lut (.A(n45730), .B(n45742), .C(n45728), 
         .D(n45735), .Z(n6_adj_509)) /* synthesis lut_function=(!(A+!((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i15777_2_lut_3_lut_4_lut_4_lut.init = 16'h5551;
    LUT4 i5478_2_lut_rep_606_4_lut_4_lut (.A(n45730), .B(n43563), .C(n895[3]), 
         .D(n2603[5]), .Z(n45727)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (D)+!B !(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5478_2_lut_rep_606_4_lut_4_lut.init = 16'h65a9;
    LUT4 div_28_i171_3_lut_4_lut (.A(n46004), .B(n22716), .C(n231[5]), 
         .D(n46022), .Z(n244)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_28_i171_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i36922_2_lut_rep_817_2_lut_3_lut_4_lut_4_lut (.A(n46001), .B(n45975), 
         .C(n45978), .D(n160), .Z(n45938)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C+(D))))) */ ;
    defparam i36922_2_lut_rep_817_2_lut_3_lut_4_lut_4_lut.init = 16'h4448;
    LUT4 i38118_2_lut_3_lut_4_lut_4_lut (.A(n46001), .B(n45953), .C(n45978), 
         .D(n160), .Z(n43883)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+!(C+(D)))) */ ;
    defparam i38118_2_lut_3_lut_4_lut_4_lut.init = 16'heeed;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_262 (.A(n45730), .B(n45724), .C(n45725), 
         .D(n45728), .Z(n43647)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_262.init = 16'hfefd;
    LUT4 i3128_3_lut_4_lut (.A(n41378), .B(n41291), .C(n45835), .D(n41360), 
         .Z(n8_adj_465)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B ((D)+!C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3128_3_lut_4_lut.init = 16'h3173;
    LUT4 i1_2_lut_2_lut_rep_822_3_lut_4_lut_4_lut (.A(n46001), .B(n45975), 
         .C(n45978), .D(n160), .Z(n45943)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+(D)))) */ ;
    defparam i1_2_lut_2_lut_rep_822_3_lut_4_lut_4_lut.init = 16'h9996;
    LUT4 i2_4_lut_adj_263 (.A(n46147), .B(n46870), .C(n31_adj_501), .D(n46589), 
         .Z(n43592)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i2_4_lut_adj_263.init = 16'h2000;
    CCU2D add_1770_5 (.A0(address[2]), .B0(n46133), .C0(n45724), .D0(akku_o_c_2), 
          .A1(address[3]), .B1(n46133), .C1(n45728), .D1(akku_o_c_3), 
          .CIN(n40406), .COUT(n40407), .S0(akku_o_8__N_50[2]), .S1(akku_o_8__N_50[3]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(79[27:57])
    defparam add_1770_5.INIT0 = 16'hd1e2;
    defparam add_1770_5.INIT1 = 16'hd1e2;
    defparam add_1770_5.INJECT1_0 = "NO";
    defparam add_1770_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_3_lut_3_lut_4_lut_4_lut (.A(n46001), .B(n45975), 
         .C(n45953), .D(n45960), .Z(n41038)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam i1_2_lut_3_lut_3_lut_3_lut_4_lut_4_lut.init = 16'h4b87;
    LUT4 i37138_1_lut_2_lut_3_lut_3_lut_3_lut_4_lut_4_lut (.A(n46001), .B(n45953), 
         .C(n45975), .D(n45960), .Z(n12)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B+!(C (D)))) */ ;
    defparam i37138_1_lut_2_lut_3_lut_3_lut_3_lut_4_lut_4_lut.init = 16'hefdf;
    LUT4 i37137_2_lut_rep_824_3_lut_4_lut_4_lut (.A(n46001), .B(n45953), 
         .C(n45975), .D(n45960), .Z(n45945)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam i37137_2_lut_rep_824_3_lut_4_lut_4_lut.init = 16'h1020;
    LUT4 i1_2_lut_rep_675_4_lut_4_lut (.A(n45888), .B(n1403[1]), .C(n45799), 
         .D(n1416[1]), .Z(n45796)) /* synthesis lut_function=(A (B (C (D))+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_rep_675_4_lut_4_lut.init = 16'ha200;
    LUT4 i1_2_lut_rep_831_3_lut_4_lut_4_lut (.A(n46001), .B(n160), .C(n45977), 
         .D(n161_adj_302), .Z(n45952)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_831_3_lut_4_lut_4_lut.init = 16'haaa9;
    LUT4 i2_3_lut_4_lut_adj_264 (.A(n45888), .B(n1403[1]), .C(n45799), 
         .D(n1416[1]), .Z(n23030)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_4_lut_adj_264.init = 16'hf708;
    LUT4 i15102_3_lut_rep_707 (.A(n45888), .B(n1403[1]), .C(n45799), .D(n1416[1]), 
         .Z(n45828)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i15102_3_lut_rep_707.init = 16'hf700;
    LUT4 div_39_i156_3_lut_rep_860_4_lut (.A(n45999), .B(n45998), .C(n45996), 
         .D(n46007), .Z(n45981)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_i156_3_lut_rep_860_4_lut.init = 16'h2fd0;
    LUT4 mux_40_i4_3_lut_rep_864_4_lut (.A(n45999), .B(n45998), .C(n11), 
         .D(n46008), .Z(n45985)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A ((D)+!C)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_40_i4_3_lut_rep_864_4_lut.init = 16'hfd0d;
    LUT4 i1_2_lut_adj_265 (.A(n39), .B(n51), .Z(n37_adj_340)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_2_lut_adj_265.init = 16'h8888;
    LUT4 i1985_2_lut (.A(address[1]), .B(address[0]), .Z(pc_5__N_35[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i1985_2_lut.init = 16'h6666;
    CCU2D add_388_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n23659), .B1(n21707), .C1(n46145), .D1(n1416[1]), .COUT(n40446), 
          .S1(n1543[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_388_1.INIT0 = 16'hF000;
    defparam add_388_1.INIT1 = 16'h07f7;
    defparam add_388_1.INJECT1_0 = "NO";
    defparam add_388_1.INJECT1_1 = "NO";
    LUT4 i23945_3_lut (.A(data[5]), .B(data[7]), .C(data[6]), .Z(n3668[1])) /* synthesis lut_function=(A ((C)+!B)+!A !(B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(90[17] 106[12])
    defparam i23945_3_lut.init = 16'hb3b3;
    LUT4 i7822_1_lut_3_lut_4_lut (.A(n45999), .B(n45998), .C(n11), .D(n46008), 
         .Z(n8_adj_464)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)))+!A ((D)+!C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i7822_1_lut_3_lut_4_lut.init = 16'h02f2;
    CCU2D add_340_7 (.A0(n1311[4]), .B0(n1311[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40445), 
          .S0(n1324[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_340_7.INIT0 = 16'h5999;
    defparam add_340_7.INIT1 = 16'h0000;
    defparam add_340_7.INJECT1_0 = "NO";
    defparam add_340_7.INJECT1_1 = "NO";
    CCU2D add_340_5 (.A0(n1311[2]), .B0(n1311[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1311[3]), .B1(n1311[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40444), .COUT(n40445), .S0(n1324[3]), .S1(n1324[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_340_5.INIT0 = 16'h5999;
    defparam add_340_5.INIT1 = 16'h5666;
    defparam add_340_5.INJECT1_0 = "NO";
    defparam add_340_5.INJECT1_1 = "NO";
    CCU2D add_1770_3 (.A0(address[0]), .B0(n46133), .C0(n45248), .D0(akku_o_c_0), 
          .A1(address[1]), .B1(n46133), .C1(n930[1]), .D1(akku_o_c_1), 
          .CIN(n40405), .COUT(n40406), .S0(n4257[0]), .S1(akku_o_8__N_50[1]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(79[27:57])
    defparam add_1770_3.INIT0 = 16'hd1e2;
    defparam add_1770_3.INIT1 = 16'hd1e2;
    defparam add_1770_3.INJECT1_0 = "NO";
    defparam add_1770_3.INJECT1_1 = "NO";
    LUT4 i37092_2_lut_rep_702_4_lut (.A(n46145), .B(n1403[1]), .C(n45888), 
         .D(n89_adj_303), .Z(n45823)) /* synthesis lut_function=(!(A ((D)+!B)+!A (((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i37092_2_lut_rep_702_4_lut.init = 16'h00c8;
    LUT4 i15850_2_lut_3_lut_4_lut (.A(n46268), .B(n46266), .C(n45_adj_356), 
         .D(n46230), .Z(n22585)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;
    defparam i15850_2_lut_3_lut_4_lut.init = 16'h0f0e;
    LUT4 i2_4_lut_4_lut_adj_266 (.A(n1403[1]), .B(n45888), .C(n45828), 
         .D(n8_adj_490), .Z(n43681)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (B (D)+!B !(C (D)+!C !(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_4_lut_4_lut_adj_266.init = 16'h12ed;
    LUT4 i3_4_lut_4_lut_adj_267 (.A(n45730), .B(n6_adj_509), .C(n2734[3]), 
         .D(n21872), .Z(n43706)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3_4_lut_4_lut_adj_267.init = 16'h9669;
    LUT4 div_53_i135_4_lut_rep_832_3_lut_4_lut (.A(n46034), .B(n46002), 
         .C(n45960), .D(n46001), .Z(n45953)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(B (C (D))+!B !(C (D))))) */ ;
    defparam div_53_i135_4_lut_rep_832_3_lut_4_lut.init = 16'h6999;
    LUT4 i1_2_lut_rep_1075_3_lut_4_lut (.A(n46264), .B(n46261), .C(n46266), 
         .D(n46268), .Z(n46196)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(39[10:22])
    defparam i1_2_lut_rep_1075_3_lut_4_lut.init = 16'hfffe;
    LUT4 i7476_2_lut_rep_856_3_lut_4_lut_4_lut (.A(n46068), .B(n46034), 
         .C(n46002), .D(n46001), .Z(n45977)) /* synthesis lut_function=(!((B (C+!(D))+!B !(C (D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i7476_2_lut_rep_856_3_lut_4_lut_4_lut.init = 16'h2800;
    LUT4 i1_2_lut_4_lut_adj_268 (.A(n1403[1]), .B(n45888), .C(n6_adj_441), 
         .D(n45828), .Z(n5_adj_507)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A !(B (C)+!B !((D)+!C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_4_lut_adj_268.init = 16'h4a7a;
    LUT4 i1_3_lut_adj_269 (.A(oprand[3]), .B(n46873), .C(oprand[2]), .Z(n4_adj_497)) /* synthesis lut_function=(!(A ((C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam i1_3_lut_adj_269.init = 16'h5d5d;
    LUT4 i31658_2_lut_rep_862_3_lut_4_lut (.A(n46006), .B(n46008), .C(n46005), 
         .D(n46007), .Z(n45983)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C+(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i31658_2_lut_rep_862_3_lut_4_lut.init = 16'hfdf0;
    LUT4 n1408_bdd_4_lut_4_lut_rep_710 (.A(n1403[1]), .B(n45888), .C(n6_adj_441), 
         .D(n45828), .Z(n45831)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B (C)+!B !(C+(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam n1408_bdd_4_lut_4_lut_rep_710.init = 16'h1f3e;
    LUT4 i2_3_lut_rep_877 (.A(n190), .B(n191), .C(n46005), .Z(n45998)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_rep_877.init = 16'hfefe;
    LUT4 i23894_2_lut_rep_871_4_lut (.A(n190), .B(n191), .C(n46005), .D(n45999), 
         .Z(n45992)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i23894_2_lut_rep_871_4_lut.init = 16'h0100;
    LUT4 rem_61_i85_3_lut_rep_1046_4_lut_4_lut_4_lut (.A(akku_o_c_3), .B(akku_o_c_2), 
         .C(akku_o_c_1), .D(akku_o_c_4), .Z(n46167)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+!(D)))+!A (B (C+!(D)))) */ ;
    defparam rem_61_i85_3_lut_rep_1046_4_lut_4_lut_4_lut.init = 16'hc2cc;
    CCU2D add_340_3 (.A0(n1311[0]), .B0(n1311[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1311[1]), .B1(n1311[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40443), .COUT(n40444), .S0(n1324[1]), .S1(n1324[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_340_3.INIT0 = 16'h5666;
    defparam add_340_3.INIT1 = 16'h5999;
    defparam add_340_3.INJECT1_0 = "NO";
    defparam add_340_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_861_3_lut_4_lut (.A(n46008), .B(n46007), .C(n46006), 
         .D(n45998), .Z(n45982)) /* synthesis lut_function=(A (B+(D))+!A !(B ((D)+!C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_rep_861_3_lut_4_lut.init = 16'haad9;
    LUT4 i1_2_lut_4_lut_adj_270 (.A(n1403[1]), .B(n45888), .C(n6_adj_441), 
         .D(n45828), .Z(n4_adj_489)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B+!(C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_4_lut_adj_270.init = 16'hefce;
    CCU2D add_340_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n43679), .B1(n7_adj_469), .C1(n46128), .D1(n510[1]), .COUT(n40443), 
          .S1(n1324[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_340_1.INIT0 = 16'hF000;
    defparam add_340_1.INIT1 = 16'h06f6;
    defparam add_340_1.INJECT1_0 = "NO";
    defparam add_340_1.INJECT1_1 = "NO";
    PFUMX i38339 (.BLUT(n45547), .ALUT(n45546), .C0(n45831), .Z(n45548));
    CCU2D add_338_7 (.A0(n1298[4]), .B0(n1298[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40442), 
          .S0(n1311[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_338_7.INIT0 = 16'h5999;
    defparam add_338_7.INIT1 = 16'h0000;
    defparam add_338_7.INJECT1_0 = "NO";
    defparam add_338_7.INJECT1_1 = "NO";
    LUT4 i15015_3_lut_4_lut (.A(n45846), .B(n45836), .C(n23490), .D(n22969), 
         .Z(n21583)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B (C+(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i15015_3_lut_4_lut.init = 16'h00ef;
    LUT4 div_46_i153_4_lut_4_lut (.A(n45997), .B(n191_adj_335), .C(n12_adj_508), 
         .D(n45984), .Z(n220_adj_405)) /* synthesis lut_function=(!(A (B+(D))+!A (B+(C+(D))))) */ ;
    defparam div_46_i153_4_lut_4_lut.init = 16'h0023;
    LUT4 i2006_2_lut_3_lut_4_lut (.A(address[2]), .B(n46277), .C(address[4]), 
         .D(address[3]), .Z(pc_5__N_35[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i2006_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 div_39_i157_3_lut_4_lut_4_lut_4_lut (.A(n46008), .B(n46007), .C(n46006), 
         .D(n45998), .Z(n224)) /* synthesis lut_function=(!(A (C)+!A !(B (C (D))+!B (C (D)+!C !(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam div_39_i157_3_lut_4_lut_4_lut_4_lut.init = 16'h5a0b;
    LUT4 i4645_2_lut_3_lut_4_lut_3_lut (.A(n720[5]), .B(n45791), .C(n46847), 
         .Z(n1947[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C)+!B !(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i4645_2_lut_3_lut_4_lut_3_lut.init = 16'hcbcb;
    LUT4 div_46_i156_3_lut_rep_852_4_lut (.A(n46042), .B(n46010), .C(n46849), 
         .D(n46009), .Z(n45973)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D)))) */ ;
    defparam div_46_i156_3_lut_rep_852_4_lut.init = 16'h9699;
    LUT4 i3_4_lut_adj_271 (.A(n122_adj_510), .B(n12888[1]), .C(n12888[2]), 
         .D(n12888[3]), .Z(n36)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i3_4_lut_adj_271.init = 16'h0002;
    LUT4 i37229_4_lut (.A(n46204), .B(n46170), .C(n46188), .D(n122_adj_510), 
         .Z(n29)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i37229_4_lut.init = 16'h0001;
    LUT4 i6621_2_lut_rep_863_3_lut_4_lut (.A(n46042), .B(n46010), .C(n45997), 
         .D(n46009), .Z(n45984)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (B (C+(D))+!B (C))) */ ;
    defparam i6621_2_lut_rep_863_3_lut_4_lut.init = 16'hf6f0;
    LUT4 pc_5__I_0_299_i1_3_lut_4_lut (.A(states[0]), .B(n46247), .C(pc[0]), 
         .D(data[0]), .Z(adress_5__N_3[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(116[33:48])
    defparam pc_5__I_0_299_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pc_5__I_0_299_i3_3_lut_4_lut (.A(states[0]), .B(n46247), .C(pc[2]), 
         .D(data[2]), .Z(adress_5__N_3[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(116[33:48])
    defparam pc_5__I_0_299_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pc_5__I_0_299_i4_3_lut_4_lut (.A(states[0]), .B(n46247), .C(pc[3]), 
         .D(data[3]), .Z(adress_5__N_3[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(116[33:48])
    defparam pc_5__I_0_299_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pc_5__I_0_299_i5_3_lut_4_lut (.A(states[0]), .B(n46247), .C(pc[4]), 
         .D(data[4]), .Z(adress_5__N_3[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(116[33:48])
    defparam pc_5__I_0_299_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pc_5__I_0_299_i6_3_lut_4_lut (.A(states[0]), .B(n46247), .C(pc[5]), 
         .D(data[5]), .Z(adress_5__N_3[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(116[33:48])
    defparam pc_5__I_0_299_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pc_5__I_0_299_i2_3_lut_4_lut (.A(states[0]), .B(n46247), .C(pc[1]), 
         .D(data[1]), .Z(adress_5__N_3[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(116[33:48])
    defparam pc_5__I_0_299_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i38149_2_lut_rep_1124 (.A(oprand[4]), .B(oprand[3]), .Z(n46245)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i38149_2_lut_rep_1124.init = 16'h7777;
    CCU2D add_1770_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n46133), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n40405));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(79[27:57])
    defparam add_1770_1.INIT0 = 16'hF000;
    defparam add_1770_1.INIT1 = 16'h0fff;
    defparam add_1770_1.INJECT1_0 = "NO";
    defparam add_1770_1.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_686_4_lut (.A(n45839), .B(n22978), .C(n43738), .D(n43762), 
         .Z(n45807)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i2_3_lut_rep_686_4_lut.init = 16'h6996;
    LUT4 i1_2_lut_rep_1089_3_lut (.A(n46873), .B(n46875), .C(n46876), 
         .Z(n46210)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_rep_1089_3_lut.init = 16'h7070;
    LUT4 i3042_4_lut_3_lut_rep_734 (.A(n43686), .B(n45856), .C(n45869), 
         .Z(n45855)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3042_4_lut_3_lut_rep_734.init = 16'h8e8e;
    LUT4 i7469_2_lut_rep_865_3_lut_4_lut (.A(n46025), .B(n130), .C(n46001), 
         .D(n46034), .Z(n45986)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i7469_2_lut_rep_865_3_lut_4_lut.init = 16'h10e0;
    LUT4 i1302_2_lut_rep_1122_3_lut (.A(\states[1] ), .B(states[0]), .C(states_c[2]), 
         .Z(n46243)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam i1302_2_lut_rep_1122_3_lut.init = 16'h0202;
    LUT4 i1298_2_lut_3_lut_4_lut (.A(\states[1] ), .B(states[0]), .C(states_c[2]), 
         .D(n4_adj_440), .Z(n3611)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam i1298_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 mux_54_i6_3_lut_4_lut (.A(n46025), .B(n130), .C(n29_adj_353), 
         .D(n46034), .Z(n218[5])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_54_i6_3_lut_4_lut.init = 16'hefe0;
    LUT4 i24151_4_lut (.A(n107), .B(n45944), .C(n270_adj_516[2]), .D(n45930), 
         .Z(n30878)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i24151_4_lut.init = 16'ha088;
    LUT4 i132_else_4_lut (.A(akku_o_c_3), .B(akku_o_c_1), .C(akku_o_c_2), 
         .Z(n46303)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i132_else_4_lut.init = 16'h0101;
    LUT4 i2_2_lut_rep_751_3_lut_4_lut_3_lut_4_lut (.A(n46019), .B(n46114), 
         .C(n45877), .D(n45924), .Z(n45872)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i2_2_lut_rep_751_3_lut_4_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i1987_2_lut_rep_1156 (.A(address[1]), .B(address[0]), .Z(n46277)) /* synthesis lut_function=(A (B)) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i1987_2_lut_rep_1156.init = 16'h8888;
    LUT4 i3513_4_lut_3_lut_4_lut (.A(n866[4]), .B(n45839), .C(n22978), 
         .D(n41108), .Z(n8_adj_420)) /* synthesis lut_function=(A (B+((D)+!C))+!A !((C+!(D))+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3513_4_lut_3_lut_4_lut.init = 16'hae8a;
    LUT4 i15392_3_lut_rep_802_4_lut (.A(n46019), .B(n46114), .C(n45924), 
         .D(n15), .Z(n45923)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;
    defparam i15392_3_lut_rep_802_4_lut.init = 16'h2220;
    LUT4 div_28_i174_3_lut_rep_859_4_lut_4_lut (.A(n217), .B(n46021), .C(n231[2]), 
         .D(n22716), .Z(n45980)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C (D))) */ ;
    defparam div_28_i174_3_lut_rep_859_4_lut_4_lut.init = 16'hf0a2;
    LUT4 div_28_i173_3_lut_4_lut_4_lut (.A(n217), .B(n46021), .C(n231[3]), 
         .D(n22716), .Z(n246_adj_458)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam div_28_i173_3_lut_4_lut_4_lut.init = 16'hf0c4;
    LUT4 mux_29_i3_3_lut_4_lut_4_lut (.A(n217), .B(n46021), .C(n7), .D(n22716), 
         .Z(n112[2])) /* synthesis lut_function=(A (B+(C+(D)))+!A !(C+!(D))) */ ;
    defparam mux_29_i3_3_lut_4_lut_4_lut.init = 16'hafa8;
    LUT4 i3114_4_lut_3_lut_rep_714 (.A(n41291), .B(n363[2]), .C(n45848), 
         .Z(n45835)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3114_4_lut_3_lut_rep_714.init = 16'h8e8e;
    LUT4 i1_2_lut_4_lut_adj_272 (.A(n46039), .B(n46030), .C(n169), .D(n190), 
         .Z(n4_adj_446)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B ((D)+!C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_4_lut_adj_272.init = 16'hffa6;
    LUT4 i1994_2_lut_rep_1116_3_lut (.A(address[1]), .B(address[0]), .C(address[2]), 
         .Z(n46237)) /* synthesis lut_function=(A (B (C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i1994_2_lut_rep_1116_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_1126 (.A(\states[1] ), .B(states_c[2]), .Z(n46247)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(116[33:48])
    defparam i1_2_lut_rep_1126.init = 16'heeee;
    LUT4 i1_2_lut_rep_1090_3_lut (.A(\states[1] ), .B(states_c[2]), .C(states[0]), 
         .Z(n46211)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(116[33:48])
    defparam i1_2_lut_rep_1090_3_lut.init = 16'hefef;
    CCU2D add_338_5 (.A0(n1298[2]), .B0(n1298[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1298[3]), .B1(n1298[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40441), .COUT(n40442), .S0(n1311[3]), .S1(n1311[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_338_5.INIT0 = 16'h5999;
    defparam add_338_5.INIT1 = 16'h5666;
    defparam add_338_5.INJECT1_0 = "NO";
    defparam add_338_5.INJECT1_1 = "NO";
    LUT4 Select_6139_i2_2_lut_rep_1054_3_lut_4_lut (.A(\states[1] ), .B(states_c[2]), 
         .C(akku_o_c_4), .D(states[0]), .Z(n46175)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(116[33:48])
    defparam Select_6139_i2_2_lut_rep_1054_3_lut_4_lut.init = 16'h1000;
    LUT4 i31638_2_lut_rep_874_3_lut (.A(n46050), .B(n169), .C(n46008), 
         .Z(n45995)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i31638_2_lut_rep_874_3_lut.init = 16'h9696;
    LUT4 rem_89_i85_3_lut_4_lut_4_lut_3_lut_4_lut (.A(akku_o_c_2), .B(akku_o_c_1), 
         .C(akku_o_c_3), .D(akku_o_c_4), .Z(n118_adj_307)) /* synthesis lut_function=(A (B+!(C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam rem_89_i85_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h8aaa;
    LUT4 i31643_2_lut_rep_875_3_lut (.A(n46050), .B(n169), .C(n46008), 
         .Z(n45996)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;
    defparam i31643_2_lut_rep_875_3_lut.init = 16'hf9f9;
    LUT4 i1_2_lut_rep_703_4_lut (.A(n41291), .B(n363[2]), .C(n45848), 
         .D(n41378), .Z(n45824)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_rep_703_4_lut.init = 16'h718e;
    LUT4 i1_2_lut_3_lut_4_lut_adj_273 (.A(n41291), .B(n363[2]), .C(n45848), 
         .D(n41378), .Z(n43727)) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_3_lut_4_lut_adj_273.init = 16'hdb24;
    LUT4 i31648_2_lut_rep_867_3_lut_4_lut_4_lut (.A(n46038), .B(n46050), 
         .C(n169), .D(n46008), .Z(n45988)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C+(D))+!B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i31648_2_lut_rep_867_3_lut_4_lut_4_lut.init = 16'h5642;
    LUT4 Select_6143_i2_2_lut_rep_1060_3_lut_4_lut (.A(\states[1] ), .B(states_c[2]), 
         .C(akku_o_c_0), .D(states[0]), .Z(n46181)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(116[33:48])
    defparam Select_6143_i2_2_lut_rep_1060_3_lut_4_lut.init = 16'h1000;
    LUT4 Select_6136_i2_2_lut_rep_1076_3_lut_4_lut (.A(\states[1] ), .B(states_c[2]), 
         .C(akku_o_c_7), .D(states[0]), .Z(n46197)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(116[33:48])
    defparam Select_6136_i2_2_lut_rep_1076_3_lut_4_lut.init = 16'h1000;
    LUT4 i3121_3_lut_rep_704_4_lut (.A(n41291), .B(n363[2]), .C(n45848), 
         .D(n41378), .Z(n45825)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (B (C (D))+!B (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3121_3_lut_rep_704_4_lut.init = 16'h04df;
    LUT4 Select_6137_i2_2_lut_rep_1077_3_lut_4_lut (.A(\states[1] ), .B(states_c[2]), 
         .C(akku_o_c_6), .D(states[0]), .Z(n46198)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(116[33:48])
    defparam Select_6137_i2_2_lut_rep_1077_3_lut_4_lut.init = 16'h1000;
    LUT4 Select_6138_i2_2_lut_rep_1078_3_lut_4_lut (.A(\states[1] ), .B(states_c[2]), 
         .C(akku_o_c_5), .D(states[0]), .Z(n46199)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(116[33:48])
    defparam Select_6138_i2_2_lut_rep_1078_3_lut_4_lut.init = 16'h1000;
    LUT4 Select_6140_i2_2_lut_rep_1079_3_lut_4_lut (.A(\states[1] ), .B(states_c[2]), 
         .C(akku_o_c_3), .D(states[0]), .Z(n46200)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(116[33:48])
    defparam Select_6140_i2_2_lut_rep_1079_3_lut_4_lut.init = 16'h1000;
    LUT4 Select_6141_i2_2_lut_rep_1080_3_lut_4_lut (.A(\states[1] ), .B(states_c[2]), 
         .C(akku_o_c_2), .D(states[0]), .Z(n46201)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(116[33:48])
    defparam Select_6141_i2_2_lut_rep_1080_3_lut_4_lut.init = 16'h1000;
    LUT4 i23760_3_lut_rep_878_4_lut_4_lut (.A(n46038), .B(n46050), .C(n169), 
         .D(n46008), .Z(n45999)) /* synthesis lut_function=(A (B+(C))+!A !(B (C+(D))+!B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i23760_3_lut_rep_878_4_lut_4_lut.init = 16'ha9bd;
    LUT4 Select_6142_i2_2_lut_rep_1081_3_lut_4_lut (.A(\states[1] ), .B(states_c[2]), 
         .C(akku_o_c_1), .D(states[0]), .Z(n46202)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(116[33:48])
    defparam Select_6142_i2_2_lut_rep_1081_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_1123_3_lut (.A(\states[1] ), .B(states_c[2]), .C(states[0]), 
         .Z(n46244)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(116[33:48])
    defparam i1_2_lut_rep_1123_3_lut.init = 16'hfefe;
    LUT4 i17177_1_lut_2_lut_3_lut (.A(\states[1] ), .B(states_c[2]), .C(states[0]), 
         .Z(clk_c_enable_26)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(116[33:48])
    defparam i17177_1_lut_2_lut_3_lut.init = 16'h0101;
    LUT4 i15488_2_lut_3_lut_4_lut (.A(\states[1] ), .B(states_c[2]), .C(n46853), 
         .D(states[0]), .Z(n22192)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(116[33:48])
    defparam i15488_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i23670_3_lut_rep_1127 (.A(akku_o_c_2), .B(akku_o_c_4), .C(akku_o_c_3), 
         .Z(n46248)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(10[13:19])
    defparam i23670_3_lut_rep_1127.init = 16'h1818;
    LUT4 i1_2_lut_rep_850_4_lut (.A(n169), .B(n46050), .C(n11), .D(n46849), 
         .Z(n45971)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A (B (D)+!B !(C (D)+!C !(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_850_4_lut.init = 16'h3ac5;
    LUT4 n6_bdd_4_lut_adj_274 (.A(n6_adj_432), .B(n2629[5]), .C(n2629[3]), 
         .D(n2629[4]), .Z(n45247)) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam n6_bdd_4_lut_adj_274.init = 16'hdb24;
    LUT4 i36945_2_lut_rep_1128 (.A(akku_o_c_1), .B(n46878), .Z(n46249)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i36945_2_lut_rep_1128.init = 16'heeee;
    LUT4 i1_2_lut_4_lut_adj_275 (.A(n41291), .B(n45848), .C(n37_adj_301), 
         .D(n23490), .Z(n41143)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_4_lut_adj_275.init = 16'h53ac;
    LUT4 i1_3_lut_4_lut_adj_276 (.A(akku_o_c_1), .B(n46878), .C(n45480), 
         .D(n31_adj_319), .Z(n43563)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_adj_276.init = 16'h1000;
    LUT4 gnd_bdd_2_lut_3_lut (.A(n46880), .B(akku_o_c_3), .C(n45721), 
         .Z(n45694)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam gnd_bdd_2_lut_3_lut.init = 16'h8080;
    LUT4 i3271_2_lut_rep_711_4_lut (.A(n41291), .B(n45848), .C(n37_adj_301), 
         .D(n45846), .Z(n45832)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B ((D)+!C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i3271_2_lut_rep_711_4_lut.init = 16'hffac;
    LUT4 i37219_2_lut_3_lut (.A(akku_o_c_3), .B(akku_o_c_0), .C(akku_o_c_2), 
         .Z(n43557)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i37219_2_lut_3_lut.init = 16'h0101;
    LUT4 i2_3_lut_3_lut_4_lut_4_lut (.A(akku_o_c_4), .B(n66), .C(akku_o_c_0), 
         .D(akku_o_c_3), .Z(n43558)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i2_3_lut_3_lut_4_lut_4_lut.init = 16'h0004;
    LUT4 i1_2_lut_rep_1129 (.A(oprand[0]), .B(oprand[3]), .Z(n46250)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_2_lut_rep_1129.init = 16'h8888;
    CCU2D add_338_3 (.A0(n1298[0]), .B0(n1298[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1298[1]), .B1(n1298[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40440), .COUT(n40441), .S0(n1311[1]), .S1(n1311[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_338_3.INIT0 = 16'h5666;
    defparam add_338_3.INIT1 = 16'h5999;
    defparam add_338_3.INJECT1_0 = "NO";
    defparam add_338_3.INJECT1_1 = "NO";
    LUT4 i6611_2_lut_rep_869_3_lut_4_lut (.A(n46031), .B(n46009), .C(n46042), 
         .Z(n45990)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i6611_2_lut_rep_869_3_lut_4_lut.init = 16'h4848;
    CCU2D add_338_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n6_adj_410), .B1(n5_adj_413), .C1(n46128), .D1(n45803), 
          .COUT(n40440), .S1(n1311[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_338_1.INIT0 = 16'hF000;
    defparam add_338_1.INIT1 = 16'h09f9;
    defparam add_338_1.INJECT1_0 = "NO";
    defparam add_338_1.INJECT1_1 = "NO";
    LUT4 i109_4_lut_3_lut (.A(oprand[0]), .B(oprand[3]), .C(oprand[4]), 
         .Z(n66)) /* synthesis lut_function=(A (B (C))+!A !(B+(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i109_4_lut_3_lut.init = 16'h8181;
    LUT4 i1_2_lut_rep_1094_3_lut (.A(n46880), .B(akku_o_c_2), .C(akku_o_c_1), 
         .Z(n46215)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_1094_3_lut.init = 16'h8080;
    FD1P3AX akku_i0_i1_rep_1179 (.D(n3555[0]), .SP(clk_c_enable_22), .CK(clk_c), 
            .Q(n46880)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam akku_i0_i1_rep_1179.GSR = "ENABLED";
    LUT4 mux_132_i6_4_lut_4_lut (.A(n45881), .B(n45840), .C(n89_adj_320), 
         .D(n545[5]), .Z(n1403[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_132_i6_4_lut_4_lut.init = 16'h8f80;
    LUT4 i1_4_lut_adj_277 (.A(n122_adj_511), .B(n117_adj_512), .C(n45404), 
         .D(n6_adj_359), .Z(n43479)) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_4_lut_adj_277.init = 16'h8020;
    LUT4 i37168_2_lut (.A(n122_adj_511), .B(n43941), .Z(n43595)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i37168_2_lut.init = 16'h1111;
    LUT4 mux_167_i6_3_lut_4_lut_4_lut_4_lut (.A(n45791), .B(n46847), .C(n19), 
         .D(n720[5]), .Z(n755[5])) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_167_i6_3_lut_4_lut_4_lut_4_lut.init = 16'hf400;
    LUT4 i23802_2_lut_3_lut_4_lut (.A(n46031), .B(n46009), .C(n46042), 
         .Z(n12_adj_508)) /* synthesis lut_function=(A ((C)+!B)+!A !(B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i23802_2_lut_3_lut_4_lut.init = 16'hb7b7;
    LUT4 i1_2_lut_rep_1035_3_lut_3_lut_4_lut_3_lut (.A(n46875), .B(n46873), 
         .C(n46876), .Z(n46156)) /* synthesis lut_function=(A (B (C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam i1_2_lut_rep_1035_3_lut_3_lut_4_lut_3_lut.init = 16'h9494;
    CCU2D add_336_7 (.A0(n1285[4]), .B0(n1285[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40439), 
          .S0(n1298[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_336_7.INIT0 = 16'h5999;
    defparam add_336_7.INIT1 = 16'h0000;
    defparam add_336_7.INJECT1_0 = "NO";
    defparam add_336_7.INJECT1_1 = "NO";
    CCU2D add_336_5 (.A0(n1285[2]), .B0(n1285[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1285[3]), .B1(n1285[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40438), .COUT(n40439), .S0(n1298[3]), .S1(n1298[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_336_5.INIT0 = 16'h5999;
    defparam add_336_5.INIT1 = 16'h5666;
    defparam add_336_5.INJECT1_0 = "NO";
    defparam add_336_5.INJECT1_1 = "NO";
    LUT4 i3499_4_lut_rep_718 (.A(n866[4]), .B(n45841), .C(n45859), .Z(n45839)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3499_4_lut_rep_718.init = 16'h8e8e;
    LUT4 rem_23_i57_3_lut_4_lut_3_lut_4_lut_3_lut (.A(n46875), .B(n46873), 
         .C(n46876), .Z(n78)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam rem_23_i57_3_lut_4_lut_3_lut_4_lut_3_lut.init = 16'h4242;
    LUT4 div_46_i155_4_lut_rep_851_3_lut_4_lut (.A(n45997), .B(n191_adj_335), 
         .C(n12_adj_508), .D(n45990), .Z(n45972)) /* synthesis lut_function=(!(A (D)+!A !(B (D)+!B (C+(D))))) */ ;
    defparam div_46_i155_4_lut_rep_851_3_lut_4_lut.init = 16'h55ba;
    LUT4 i1_2_lut_rep_712_4_lut (.A(n866[4]), .B(n45841), .C(n45859), 
         .D(n22978), .Z(n45833)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_rep_712_4_lut.init = 16'h718e;
    LUT4 div_46_i154_3_lut_4_lut_4_lut (.A(n45997), .B(n191_adj_335), .C(n12_adj_508), 
         .D(n45990), .Z(n221_adj_435)) /* synthesis lut_function=(A (B)+!A (B (D)+!B !(C+(D)))) */ ;
    defparam div_46_i154_3_lut_4_lut_4_lut.init = 16'hcc89;
    LUT4 mux_47_i5_3_lut_rep_880_4_lut (.A(n46031), .B(n46123), .C(n46009), 
         .Z(n46001)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_47_i5_3_lut_rep_880_4_lut.init = 16'he2e2;
    LUT4 i2_2_lut (.A(n6_adj_341), .B(n2203[5]), .Z(n7_adj_392)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i2_2_lut.init = 16'h6666;
    LUT4 i24325_2_lut_rep_1072_3_lut_4_lut (.A(oprand[1]), .B(oprand[2]), 
         .C(oprand[4]), .D(oprand[3]), .Z(n46193)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i24325_2_lut_rep_1072_3_lut_4_lut.init = 16'hf080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_278 (.A(oprand[1]), .B(oprand[2]), .C(oprand[3]), 
         .D(oprand[4]), .Z(n117_adj_512)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A !((D)+!C)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_278.init = 16'h80f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_279 (.A(oprand[1]), .B(oprand[2]), .C(oprand[3]), 
         .D(oprand[4]), .Z(n77)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (C+!(D))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_279.init = 16'hf8ff;
    LUT4 i1_2_lut_3_lut_4_lut_adj_280 (.A(oprand[1]), .B(oprand[2]), .C(oprand[4]), 
         .D(oprand[3]), .Z(n30168)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (C+!(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_280.init = 16'h0700;
    LUT4 i3506_4_lut_rep_713_4_lut (.A(n866[4]), .B(n45841), .C(n45859), 
         .D(n22978), .Z(n45834)) /* synthesis lut_function=(A (B+!(C (D)))+!A !((C+(D))+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3506_4_lut_rep_713_4_lut.init = 16'h8aae;
    LUT4 i1_2_lut_rep_1135 (.A(n46876), .B(n46875), .Z(n46256)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam i1_2_lut_rep_1135.init = 16'h8888;
    LUT4 mux_146_i4_3_lut_rep_669 (.A(n1556[5]), .B(n615[3]), .C(n89_adj_303), 
         .Z(n45790)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_146_i4_3_lut_rep_669.init = 16'h5c5c;
    LUT4 i170_2_lut_rep_1065_3_lut_4_lut (.A(oprand[2]), .B(oprand[3]), 
         .C(oprand[1]), .D(oprand[4]), .Z(n46186)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam i170_2_lut_rep_1065_3_lut_4_lut.init = 16'h0700;
    LUT4 i1_2_lut_rep_1088_3_lut (.A(oprand[2]), .B(oprand[3]), .C(oprand[4]), 
         .Z(n46209)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam i1_2_lut_rep_1088_3_lut.init = 16'h7070;
    LUT4 mux_72_i6_3_lut_rep_819_4_lut (.A(n46081), .B(n46019), .C(n43592), 
         .D(n293[1]), .Z(n45940)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam mux_72_i6_3_lut_rep_819_4_lut.init = 16'h8f80;
    LUT4 i1999_2_lut_3_lut_4_lut (.A(address[1]), .B(address[0]), .C(address[3]), 
         .D(address[2]), .Z(pc_5__N_35[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i1999_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_281 (.A(n866[4]), .B(n45841), .C(n45859), 
         .D(n22978), .Z(n41285)) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_3_lut_4_lut_adj_281.init = 16'hdb24;
    LUT4 i5463_2_lut_rep_612_3_lut_3_lut (.A(n45771), .B(n45749), .C(n46845), 
         .Z(n45733)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5463_2_lut_rep_612_3_lut_3_lut.init = 16'hf7f7;
    LUT4 i2_3_lut_4_lut_adj_282 (.A(n46081), .B(n46019), .C(n45915), .D(n293[1]), 
         .Z(n22852)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_4_lut_adj_282.init = 16'hf708;
    LUT4 i14959_3_lut_4_lut_rep_892 (.A(n46081), .B(n46019), .C(n45915), 
         .D(n293[1]), .Z(n46013)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i14959_3_lut_4_lut_rep_892.init = 16'hf700;
    CCU2D add_336_3 (.A0(n1285[0]), .B0(n1285[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1285[1]), .B1(n1285[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40437), .COUT(n40438), .S0(n1298[1]), .S1(n1298[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_336_3.INIT0 = 16'h5666;
    defparam add_336_3.INIT1 = 16'h5999;
    defparam add_336_3.INJECT1_0 = "NO";
    defparam add_336_3.INJECT1_1 = "NO";
    LUT4 i4051_2_lut_rep_717_4_lut (.A(n4_adj_389), .B(n45883), .C(n4217[1]), 
         .D(n45881), .Z(n45838)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i4051_2_lut_rep_717_4_lut.init = 16'h20ff;
    LUT4 i2_3_lut_rep_787_4_lut (.A(n46081), .B(n46019), .C(n45915), .D(n293[1]), 
         .Z(n45908)) /* synthesis lut_function=(!(A (B (C (D))+!B (D))+!A !(B+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_rep_787_4_lut.init = 16'h5dee;
    LUT4 i24311_2_lut_rep_1067_3_lut_4_lut (.A(oprand[2]), .B(oprand[3]), 
         .C(oprand[1]), .D(oprand[4]), .Z(n46188)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam i24311_2_lut_rep_1067_3_lut_4_lut.init = 16'h70f0;
    LUT4 oprand_2__bdd_3_lut_rep_1083_4_lut_4_lut (.A(oprand[2]), .B(oprand[3]), 
         .C(n46878), .D(oprand[4]), .Z(n46204)) /* synthesis lut_function=(!((B (C (D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam oprand_2__bdd_3_lut_rep_1083_4_lut_4_lut.init = 16'h2aaa;
    LUT4 i1_2_lut_rep_815_4_lut_4_lut (.A(n46019), .B(n43592), .C(n293[1]), 
         .D(n46012), .Z(n45936)) /* synthesis lut_function=(A (B (D)+!B !(C))+!A (B (D)+!B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_815_4_lut_4_lut.init = 16'hde12;
    LUT4 i1_2_lut_rep_1136 (.A(oprand[2]), .B(oprand[3]), .C(oprand[4]), 
         .Z(n46257)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam i1_2_lut_rep_1136.init = 16'h8080;
    LUT4 mux_100_i5_3_lut_rep_720 (.A(n23490), .B(n45849), .C(n15_adj_316), 
         .Z(n45841)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_100_i5_3_lut_rep_720.init = 16'hc5c5;
    LUT4 i1_2_lut_3_lut_4_lut_adj_283 (.A(n46019), .B(n43592), .C(n4201[1]), 
         .D(n45940), .Z(n405[2])) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_3_lut_4_lut_adj_283.init = 16'h0f2d;
    LUT4 i4417_2_lut_rep_663_4_lut (.A(n1556[5]), .B(n615[3]), .C(n89_adj_303), 
         .D(n1687[5]), .Z(n45784)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(B (D)+!B (C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i4417_2_lut_rep_663_4_lut.init = 16'ha35c;
    LUT4 rem_101_i84_3_lut_rep_1049_4_lut_4_lut_4_lut (.A(oprand[2]), .B(oprand[3]), 
         .C(oprand[4]), .D(oprand[1]), .Z(n46170)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:22])
    defparam rem_101_i84_3_lut_rep_1049_4_lut_4_lut_4_lut.init = 16'h4ccc;
    LUT4 n264_bdd_4_lut_38297 (.A(n261[6]), .B(n261[5]), .C(n261[8]), 
         .D(n261[4]), .Z(n45461)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n264_bdd_4_lut_38297.init = 16'hfffe;
    LUT4 i5647_4_lut_4_lut (.A(n2098[1]), .B(n2098[5]), .C(n2098[0]), 
         .D(n755[0]), .Z(n4_adj_347)) /* synthesis lut_function=(A ((C (D))+!B)+!A !(B+!(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5647_4_lut_4_lut.init = 16'hb332;
    LUT4 i15624_2_lut_rep_1137 (.A(akku_o_c_3), .B(akku_o_c_4), .Z(n46258)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i15624_2_lut_rep_1137.init = 16'h8888;
    LUT4 i14929_2_lut_rep_812_3_lut_4_lut (.A(n46019), .B(n43592), .C(n4201[1]), 
         .D(n45940), .Z(n45933)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i14929_2_lut_rep_812_3_lut_4_lut.init = 16'hf0d0;
    LUT4 i2539_2_lut_rep_814_4_lut_3_lut (.A(n46019), .B(n43592), .C(n293[1]), 
         .Z(n45935)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i2539_2_lut_rep_814_4_lut_3_lut.init = 16'hfdfd;
    LUT4 i15785_2_lut_rep_1085_3_lut (.A(akku_o_c_3), .B(akku_o_c_4), .C(akku_o_c_2), 
         .Z(n46206)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i15785_2_lut_rep_1085_3_lut.init = 16'h7070;
    CCU2D add_336_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n46870), .B1(n45804), .C1(n43341), .D1(n45806), .COUT(n40437), 
          .S1(n1298[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_336_1.INIT0 = 16'hF000;
    defparam add_336_1.INIT1 = 16'h04fe;
    defparam add_336_1.INJECT1_0 = "NO";
    defparam add_336_1.INJECT1_1 = "NO";
    LUT4 mux_160_i5_3_lut_rep_670 (.A(n1816[5]), .B(n685[4]), .C(n89), 
         .Z(n45791)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_160_i5_3_lut_rep_670.init = 16'h5c5c;
    LUT4 mux_93_i2_3_lut_4_lut (.A(n45845), .B(n15), .C(n37_adj_301), 
         .D(n45810), .Z(n396[1])) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_93_i2_3_lut_4_lut.init = 16'h08f8;
    LUT4 i5848_2_lut_3_lut_4_lut (.A(n45845), .B(n15), .C(n363[0]), .D(n45810), 
         .Z(n9959)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i5848_2_lut_3_lut_4_lut.init = 16'h7000;
    LUT4 i5849_2_lut_3_lut_4_lut (.A(n45845), .B(n15), .C(n363[0]), .D(n45810), 
         .Z(n21937)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i5849_2_lut_3_lut_4_lut.init = 16'hfff7;
    LUT4 i15156_3_lut_4_lut (.A(n46026), .B(n46040), .C(n46138), .D(n43564), 
         .Z(n2293[1])) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (((D)+!C)+!B))) */ ;
    defparam i15156_3_lut_4_lut.init = 16'h0060;
    CCU2D add_334_7 (.A0(n40857), .B0(n545[8]), .C0(n45886), .D0(n45840), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40436), 
          .S0(n1285[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_334_7.INIT0 = 16'ha955;
    defparam add_334_7.INIT1 = 16'h0000;
    defparam add_334_7.INJECT1_0 = "NO";
    defparam add_334_7.INJECT1_1 = "NO";
    LUT4 i2_3_lut_4_lut_adj_284 (.A(n45753), .B(n45750), .C(n790[2]), 
         .D(n2216[2]), .Z(n40766)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A !(B (D)+!B !(C (D)+!C !(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_4_lut_adj_284.init = 16'h6798;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_285 (.A(n46033), .B(n825[7]), .C(n2293[1]), 
         .D(n45781), .Z(n23068)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A !(B (C (D))+!B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_285.init = 16'h8747;
    CCU2D add_334_5 (.A0(n45653), .B0(n45886), .C0(n545[8]), .D0(n45840), 
          .A1(n45881), .B1(n45838), .C1(n45883), .D1(n45652), .CIN(n40435), 
          .COUT(n40436), .S0(n1285[3]), .S1(n1285[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_334_5.INIT0 = 16'h56aa;
    defparam add_334_5.INIT1 = 16'h9669;
    defparam add_334_5.INJECT1_0 = "NO";
    defparam add_334_5.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_689_4_lut (.A(n45847), .B(n640[1]), .C(n43732), 
         .D(n43765), .Z(n45810)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i2_3_lut_rep_689_4_lut.init = 16'h6996;
    LUT4 oprand_3__bdd_3_lut_38564 (.A(oprand[2]), .B(oprand[0]), .C(oprand[4]), 
         .Z(n45479)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam oprand_3__bdd_3_lut_38564.init = 16'h0101;
    LUT4 i5075_2_lut_3_lut_4_lut_4_lut (.A(n46033), .B(n825[7]), .C(n2293[1]), 
         .D(n45781), .Z(n8_adj_442)) /* synthesis lut_function=(((C (D))+!B)+!A) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i5075_2_lut_3_lut_4_lut_4_lut.init = 16'hf777;
    LUT4 i1_3_lut_4_lut_adj_286 (.A(akku_o_c_2), .B(akku_o_c_1), .C(akku_o_c_4), 
         .D(akku_o_c_3), .Z(n117_adj_305)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i1_3_lut_4_lut_adj_286.init = 16'h1f00;
    LUT4 i1_3_lut_4_lut_adj_287 (.A(akku_o_c_2), .B(akku_o_c_1), .C(akku_o_c_3), 
         .D(akku_o_c_4), .Z(n5)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i1_3_lut_4_lut_adj_287.init = 16'h1f00;
    LUT4 i3092_3_lut_4_lut (.A(n640[1]), .B(n45850), .C(n45847), .D(n640[2]), 
         .Z(n8_adj_423)) /* synthesis lut_function=(A ((C (D))+!B)+!A !(B+!(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3092_3_lut_4_lut.init = 16'hb332;
    LUT4 i7486_2_lut_rep_857_4_lut_then_4_lut (.A(n46001), .B(n46034), .C(n130), 
         .D(n46850), .Z(n46307)) /* synthesis lut_function=(!(A (B (D)+!B !(C+(D)))+!A (B ((D)+!C)+!B !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i7486_2_lut_rep_857_4_lut_then_4_lut.init = 16'h33e8;
    LUT4 i33700_2_lut_rep_1070_3_lut_4_lut_4_lut (.A(akku_o_c_2), .B(akku_o_c_1), 
         .C(akku_o_c_4), .D(akku_o_c_3), .Z(n46191)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A ((C (D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i33700_2_lut_rep_1070_3_lut_4_lut_4_lut.init = 16'h2ccc;
    LUT4 mux_1263_i7_4_lut (.A(n22207), .B(akku_o_8__N_67[6]), .C(n46243), 
         .D(n3611), .Z(n3555[6])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(73[13] 82[22])
    defparam mux_1263_i7_4_lut.init = 16'hc0ca;
    LUT4 i24002_2_lut_rep_1043_3_lut_4_lut_4_lut (.A(akku_o_c_2), .B(akku_o_c_1), 
         .C(akku_o_c_0), .D(n46258), .Z(n46164)) /* synthesis lut_function=(A (B (C+!(D))+!B (C+(D)))+!A (B (C+!(D))+!B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[39:53])
    defparam i24002_2_lut_rep_1043_3_lut_4_lut_4_lut.init = 16'hf2fc;
    LUT4 i1_4_lut_adj_288 (.A(n122), .B(n46173), .C(n46358), .D(akku_o_c_0), 
         .Z(n43481)) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[8:32])
    defparam i1_4_lut_adj_288.init = 16'h8020;
    LUT4 i15503_4_lut (.A(akku_o_c_6), .B(akku_o_8__N_50[6]), .C(states_c[2]), 
         .D(data[6]), .Z(n22207)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(73[13] 82[22])
    defparam i15503_4_lut.init = 16'hc0c5;
    LUT4 i23854_2_lut_rep_721_4_lut (.A(n449[4]), .B(n3[1]), .C(n37_adj_340), 
         .D(n15), .Z(n45842)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (D)+!B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i23854_2_lut_rep_721_4_lut.init = 16'h5c00;
    LUT4 i33698_2_lut_rep_1042_3_lut_3_lut_4_lut_4_lut (.A(oprand[1]), .B(oprand[2]), 
         .C(oprand[3]), .D(oprand[4]), .Z(n46163)) /* synthesis lut_function=(!(A (C (D))+!A !(B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(20[15:21])
    defparam i33698_2_lut_rep_1042_3_lut_3_lut_4_lut_4_lut.init = 16'h4aaa;
    CCU2D add_334_3 (.A0(n45881), .B0(n45838), .C0(n545[5]), .D0(GND_net), 
          .A1(n21696), .B1(n45886), .C1(n545[8]), .D1(n45840), .CIN(n40434), 
          .COUT(n40435), .S0(n1285[1]), .S1(n1285[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_334_3.INIT0 = 16'h9969;
    defparam add_334_3.INIT1 = 16'h56aa;
    defparam add_334_3.INJECT1_0 = "NO";
    defparam add_334_3.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_adj_289 (.A(n46878), .B(oprand[2]), .C(oprand[3]), 
         .D(oprand[4]), .Z(n10)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(20[15:21])
    defparam i1_3_lut_4_lut_adj_289.init = 16'h1f00;
    LUT4 mux_1263_i8_4_lut (.A(n22209), .B(akku_o_8__N_67[7]), .C(n46243), 
         .D(n3611), .Z(n3555[7])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(73[13] 82[22])
    defparam mux_1263_i8_4_lut.init = 16'hc0ca;
    LUT4 i1_3_lut_4_lut_adj_290 (.A(oprand[1]), .B(oprand[2]), .C(oprand[4]), 
         .D(n46875), .Z(n117)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(20[15:21])
    defparam i1_3_lut_4_lut_adj_290.init = 16'h1f00;
    LUT4 i38124_2_lut_rep_1002_4_lut_then_3_lut_4_lut (.A(oprand[0]), .B(akku_o_c_0), 
         .C(oprand[1]), .D(n43), .Z(n46861)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i38124_2_lut_rep_1002_4_lut_then_3_lut_4_lut.init = 16'hefff;
    LUT4 i5427_2_lut_rep_624_3_lut_3_lut_4_lut (.A(n43563), .B(n46130), 
         .C(n45749), .D(n45771), .Z(n45745)) /* synthesis lut_function=(A (C+!(D))+!A (B+(C+!(D)))) */ ;
    defparam i5427_2_lut_rep_624_3_lut_3_lut_4_lut.init = 16'hf4ff;
    LUT4 i5381_2_lut_rep_647_4_lut_4_lut (.A(n43563), .B(n46130), .C(n45778), 
         .D(n45773), .Z(n45768)) /* synthesis lut_function=(!(A (D)+!A !(B+(C)))) */ ;
    defparam i5381_2_lut_rep_647_4_lut_4_lut.init = 16'h54fe;
    LUT4 i24314_2_lut_rep_1140 (.A(n46876), .B(n46875), .Z(n46261)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24314_2_lut_rep_1140.init = 16'heeee;
    LUT4 i38085_2_lut_3_lut_4_lut_4_lut_3_lut_4_lut (.A(n43563), .B(n46130), 
         .C(n45749), .D(n45771), .Z(n44713)) /* synthesis lut_function=(!(A (C (D))+!A (B+(C (D))))) */ ;
    defparam i38085_2_lut_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h0bbb;
    LUT4 i15505_4_lut (.A(akku_o_c_7), .B(akku_o_8__N_50[7]), .C(states_c[2]), 
         .D(data[7]), .Z(n22209)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(73[13] 82[22])
    defparam i15505_4_lut.init = 16'hc0c5;
    LUT4 i2_3_lut_4_lut_adj_291 (.A(n449[4]), .B(n3[0]), .C(n3[1]), .D(n41411), 
         .Z(n42171)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_4_lut_adj_291.init = 16'h8a00;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_adj_292 (.A(n43563), .B(n46130), .C(n45749), 
         .D(n45771), .Z(n23553)) /* synthesis lut_function=(!(A (C (D))+!A !(B (C (D))+!B !(C (D))))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut_adj_292.init = 16'h4bbb;
    LUT4 i37189_3_lut_4_lut (.A(n449[4]), .B(n3[0]), .C(n3[1]), .D(n41411), 
         .Z(n44079)) /* synthesis lut_function=(A+(B ((D)+!C)+!B (D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i37189_3_lut_4_lut.init = 16'hffae;
    LUT4 i3266_3_lut_4_lut (.A(n45849), .B(n45861), .C(n45836), .D(n23490), 
         .Z(n776[2])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i3266_3_lut_4_lut.init = 16'h6966;
    LUT4 i15144_4_lut_4_lut_rep_644_3_lut (.A(n45789), .B(n45787), .C(n45761), 
         .Z(n45765)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i15144_4_lut_4_lut_rep_644_3_lut.init = 16'h6060;
    LUT4 i1_3_lut_rep_1091_3_lut (.A(n46876), .B(oprand[3]), .C(oprand[4]), 
         .Z(n46212)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;
    defparam i1_3_lut_rep_1091_3_lut.init = 16'h4a4a;
    LUT4 mux_1263_i9_4_lut (.A(n22210), .B(akku_o_8__N_67[8]), .C(n46243), 
         .D(n3611), .Z(n3555[8])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(73[13] 82[22])
    defparam mux_1263_i9_4_lut.init = 16'hc0ca;
    LUT4 i1_4_lut_4_lut_4_lut_3_lut (.A(oprand[2]), .B(n46875), .C(oprand[4]), 
         .Z(n9_adj_487)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_4_lut_4_lut_4_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_4_lut_4_lut_adj_293 (.A(oprand[2]), .B(oprand[3]), .C(oprand[1]), 
         .D(oprand[4]), .Z(n4_adj_500)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B (C (D))))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_293.init = 16'h40a0;
    LUT4 i15506_4_lut (.A(akku_o_8__N_50[8]), .B(n895[8]), .C(n46133), 
         .D(n4_adj_513), .Z(n22210)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(73[13] 82[22])
    defparam i15506_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut_adj_294 (.A(n43563), .B(\states[1] ), .Z(n4_adj_513)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_adj_294.init = 16'h4444;
    LUT4 i33678_2_lut_rep_1045_3_lut_3_lut_4_lut (.A(n46876), .B(oprand[3]), 
         .C(n46873), .D(oprand[1]), .Z(n46166)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;
    defparam i33678_2_lut_rep_1045_3_lut_3_lut_4_lut.init = 16'h0fe0;
    LUT4 i24345_2_lut_rep_1074_3_lut_4_lut (.A(oprand[2]), .B(n46875), .C(oprand[0]), 
         .D(n46878), .Z(n46195)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24345_2_lut_rep_1074_3_lut_4_lut.init = 16'hfffe;
    LUT4 i37282_2_lut (.A(n122), .B(n44162), .Z(n43598)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i37282_2_lut.init = 16'h1111;
    LUT4 i23853_2_lut_rep_893_4_lut (.A(n46027), .B(n46056), .C(n37_adj_318), 
         .D(n43592), .Z(n46014)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B (D)+!B ((D)+!C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i23853_2_lut_rep_893_4_lut.init = 16'h005c;
    LUT4 i1_2_lut_rep_882_4_lut (.A(n46027), .B(n46056), .C(n37_adj_318), 
         .D(n46114), .Z(n46003)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B (D)+!B ((D)+!C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_882_4_lut.init = 16'h005c;
    LUT4 i2378_2_lut_rep_891_4_lut (.A(n46027), .B(n46056), .C(n37_adj_318), 
         .D(n46081), .Z(n46012)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (D)+!B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i2378_2_lut_rep_891_4_lut.init = 16'h5c00;
    PFUMX i38513 (.BLUT(n46407), .ALUT(n46408), .C0(n46014), .Z(n46409));
    LUT4 i15812_4_lut (.A(akku_o_c_1), .B(akku_o_8__N_67[1]), .C(n46276), 
         .D(data[1]), .Z(n22539)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(73[13] 82[22])
    defparam i15812_4_lut.init = 16'hc0c5;
    LUT4 i1_2_lut_3_lut_adj_295 (.A(address[1]), .B(address[0]), .C(address[2]), 
         .Z(n23757)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i1_2_lut_3_lut_adj_295.init = 16'hf7f7;
    PFUMX i38511 (.BLUT(n46404), .ALUT(n46405), .C0(n1582[3]), .Z(n46406));
    LUT4 i1_2_lut_rep_798_3_lut_4_lut (.A(n23063), .B(n46046), .C(n43683), 
         .D(n4_adj_317), .Z(n45919)) /* synthesis lut_function=(!(A (C)+!A !(B (C (D)+!C !(D))+!B !(C)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i1_2_lut_rep_798_3_lut_4_lut.init = 16'h4b0f;
    LUT4 i15111_4_lut (.A(n46043), .B(n46137), .C(n46051), .D(n46115), 
         .Z(n4382[1])) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i15111_4_lut.init = 16'h4888;
    PFUMX i38509 (.BLUT(n46245), .ALUT(n46402), .C0(n46882), .Z(n46403));
    LUT4 i1992_2_lut_3_lut (.A(address[1]), .B(address[0]), .C(address[2]), 
         .Z(pc_5__N_35[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // C:/lscc/diamond/3.11_x64/ispfpga/vhdl_packages/numeric_std.vhd(1241[12:13])
    defparam i1992_2_lut_3_lut.init = 16'h7878;
    PFUMX i38507 (.BLUT(n46398), .ALUT(n46399), .C0(n1051[3]), .Z(n46400));
    PFUMX i38505 (.BLUT(n46395), .ALUT(n46396), .C0(n208[1]), .Z(n46397));
    LUT4 div_39_i135_3_lut_rep_886_4_lut (.A(n46078), .B(n46053), .C(n169), 
         .D(n46050), .Z(n46007)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+(D))))) */ ;
    defparam div_39_i135_3_lut_rep_886_4_lut.init = 16'h6669;
    LUT4 i24251_2_lut_rep_908_3_lut_4_lut (.A(n46143), .B(n46852), .C(n22715), 
         .D(n46155), .Z(n46029)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C))+!A (B (C)+!B (C+(D))))) */ ;
    defparam i24251_2_lut_rep_908_3_lut_4_lut.init = 16'h060f;
    PFUMX i38501 (.BLUT(n46389), .ALUT(n46390), .C0(oprand[4]), .Z(n45287));
    LUT4 i6468_2_lut_rep_902_3_lut_4_lut_4_lut (.A(n46089), .B(n46078), 
         .C(n46053), .D(n46050), .Z(n46023)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+!(D)))+!A !(B+!(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i6468_2_lut_rep_902_3_lut_4_lut_4_lut.init = 16'h9a18;
    PFUMX i38499 (.BLUT(n46386), .ALUT(n46387), .C0(n46266), .Z(n46388));
    LUT4 i15806_4_lut (.A(akku_o_8__N_50[3]), .B(n45725), .C(n46854), 
         .D(n3622), .Z(n22533)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(73[13] 82[22])
    defparam i15806_4_lut.init = 16'hca0a;
    LUT4 i2_3_lut_4_lut_4_lut_adj_296 (.A(n3[3]), .B(n45866), .C(n3[2]), 
         .D(n427[1]), .Z(n41077)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2_3_lut_4_lut_4_lut_adj_296.init = 16'he718;
    PFUMX i38497 (.BLUT(n46383), .ALUT(n46384), .C0(n46876), .Z(n46385));
    LUT4 i15816_4_lut (.A(akku_o_c_3), .B(akku_o_8__N_67[3]), .C(n46276), 
         .D(data[3]), .Z(n22543)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(73[13] 82[22])
    defparam i15816_4_lut.init = 16'hc0c5;
    PFUMX i38495 (.BLUT(n46380), .ALUT(n46381), .C0(n45951), .Z(n46382));
    LUT4 i15804_4_lut (.A(akku_o_8__N_50[2]), .B(n43708), .C(n46854), 
         .D(n3622), .Z(n22531)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(73[13] 82[22])
    defparam i15804_4_lut.init = 16'hca0a;
    LUT4 i1_4_lut_4_lut_adj_297 (.A(oprand[3]), .B(oprand[4]), .C(oprand[2]), 
         .D(oprand[1]), .Z(n30180)) /* synthesis lut_function=(A (B (C (D))+!B !(C+!(D)))+!A !(B+!(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(20[15:21])
    defparam i1_4_lut_4_lut_adj_297.init = 16'h9300;
    PFUMX i38493 (.BLUT(n46309), .ALUT(n46378), .C0(akku_o_c_4), .Z(n46379));
    LUT4 mux_86_i5_3_lut_rep_735 (.A(n541[4]), .B(n45877), .C(n15), .Z(n45856)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam mux_86_i5_3_lut_rep_735.init = 16'hc5c5;
    FD1P3AX oprand_i0_i1_rep_1177 (.D(data[1]), .SP(clk_c_enable_26), .CK(clk_c), 
            .Q(n46878)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam oprand_i0_i1_rep_1177.GSR = "ENABLED";
    PFUMX i38491 (.BLUT(n46383), .ALUT(n46375), .C0(n46876), .Z(n46376));
    LUT4 i38268_then_3_lut (.A(akku_o_c_3), .B(akku_o_c_2), .C(akku_o_c_1), 
         .Z(n46310)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i38268_then_3_lut.init = 16'h0101;
    PFUMX i38489 (.BLUT(n46371), .ALUT(n46372), .C0(n45889), .Z(n1687[5]));
    LUT4 i37180_3_lut_4_lut (.A(n46051), .B(n46104), .C(n755[6]), .D(n43564), 
         .Z(n23051)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((D)+!C))) */ ;
    defparam i37180_3_lut_4_lut.init = 16'h0078;
    PFUMX i38487 (.BLUT(n46368), .ALUT(n46369), .C0(n46873), .Z(n46370));
    LUT4 i38268_else_3_lut (.A(akku_o_c_3), .B(akku_o_c_2), .C(n46880), 
         .D(akku_o_c_1), .Z(n46309)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i38268_else_3_lut.init = 16'h0001;
    PFUMX i38485 (.BLUT(n46365), .ALUT(n46366), .C0(akku_o_c_1), .Z(n46367));
    LUT4 i37044_1_lut_2_lut_3_lut_4_lut (.A(n46051), .B(n46104), .C(n46041), 
         .D(n46090), .Z(n8_adj_477)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (C (D)))) */ ;
    defparam i37044_1_lut_2_lut_3_lut_4_lut.init = 16'h0777;
    PFUMX i38483 (.BLUT(n46362), .ALUT(n46363), .C0(n43564), .Z(n46364));
    PFUMX i38481 (.BLUT(n46359), .ALUT(n46360), .C0(n790[2]), .Z(n6_adj_341));
    LUT4 i37043_2_lut_rep_894_3_lut_4_lut (.A(n46051), .B(n46104), .C(n46041), 
         .D(n46090), .Z(n46015)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;
    defparam i37043_2_lut_rep_894_3_lut_4_lut.init = 16'hf888;
    PFUMX i38479 (.BLUT(n46356), .ALUT(n46357), .C0(akku_o_c_0), .Z(n46358));
    CCU2D add_334_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n45896), .B1(n46051), .C1(n46128), .D1(n1156[1]), .COUT(n40434), 
          .S1(n1285[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_334_1.INIT0 = 16'hF000;
    defparam add_334_1.INIT1 = 16'h07f7;
    defparam add_334_1.INJECT1_0 = "NO";
    defparam add_334_1.INJECT1_1 = "NO";
    CCU2D add_283_7 (.A0(n1038[4]), .B0(n1038[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40433), 
          .S0(n1051[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_283_7.INIT0 = 16'h5999;
    defparam add_283_7.INIT1 = 16'h0000;
    defparam add_283_7.INJECT1_0 = "NO";
    defparam add_283_7.INJECT1_1 = "NO";
    PFUMX i38477 (.BLUT(n46353), .ALUT(n46354), .C0(akku_o_c_3), .Z(n45390));
    PFUMX i38475 (.BLUT(n46350), .ALUT(n46351), .C0(oprand[1]), .Z(n6_adj_359));
    LUT4 i24249_4_lut (.A(n46124), .B(n46145), .C(n46051), .D(n45896), 
         .Z(n4_adj_403)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i24249_4_lut.init = 16'h8880;
    LUT4 i1_2_lut_rep_905_4_lut (.A(n43547), .B(n46052), .C(n46137), .D(n46090), 
         .Z(n46026)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i1_2_lut_rep_905_4_lut.init = 16'h8000;
    LUT4 i2_3_lut_4_lut_adj_298 (.A(n46052), .B(n46090), .C(n46044), .D(n46137), 
         .Z(n4382[2])) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i2_3_lut_4_lut_adj_298.init = 16'h8000;
    LUT4 mux_22_i6_3_lut_4_lut (.A(oprand[0]), .B(akku_o_c_0), .C(n16[6]), 
         .D(n16[5]), .Z(n124)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_22_i6_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_2_lut_rep_1003_3_lut_4_lut (.A(n46882), .B(n46880), .C(n89_adj_320), 
         .D(n43341), .Z(n46124)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;
    defparam i1_2_lut_rep_1003_3_lut_4_lut.init = 16'h0f0e;
    PFUMX i38471 (.BLUT(n46343), .ALUT(n46344), .C0(n46878), .Z(n46345));
    LUT4 i15814_4_lut (.A(akku_o_c_2), .B(akku_o_8__N_67[2]), .C(n46276), 
         .D(data[2]), .Z(n22541)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(73[13] 82[22])
    defparam i15814_4_lut.init = 16'hc0c5;
    CCU2D add_283_5 (.A0(n1038[2]), .B0(n1038[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1038[3]), .B1(n1038[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40432), .COUT(n40433), .S0(n1051[3]), .S1(n1051[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_283_5.INIT0 = 16'h5999;
    defparam add_283_5.INIT1 = 16'h5666;
    defparam add_283_5.INJECT1_0 = "NO";
    defparam add_283_5.INJECT1_1 = "NO";
    CCU2D add_283_3 (.A0(n1038[0]), .B0(n1038[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1038[1]), .B1(n1038[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40431), .COUT(n40432), .S0(n1051[1]), .S1(n1051[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_283_3.INIT0 = 16'h5999;
    defparam add_283_3.INIT1 = 16'h5999;
    defparam add_283_3.INJECT1_0 = "NO";
    defparam add_283_3.INJECT1_1 = "NO";
    PFUMX i38469 (.BLUT(n46340), .ALUT(n46341), .C0(oprand[4]), .Z(n46342));
    LUT4 i23884_2_lut_rep_999_3_lut (.A(n46882), .B(n46880), .C(n7), .Z(n46120)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i23884_2_lut_rep_999_3_lut.init = 16'he0e0;
    PFUMX i38467 (.BLUT(n46337), .ALUT(n46338), .C0(n46875), .Z(n46339));
    LUT4 i1_2_lut_rep_1017_3_lut_4_lut (.A(n46882), .B(n46880), .C(n43668), 
         .D(n43655), .Z(n46138)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_1017_3_lut_4_lut.init = 16'hfffe;
    CCU2D add_283_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n46229), .B1(n46230), .C1(n462[1]), .D1(n462[5]), .COUT(n40431), 
          .S1(n1051[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_283_1.INIT0 = 16'hF000;
    defparam add_283_1.INIT1 = 16'h0e1f;
    defparam add_283_1.INJECT1_0 = "NO";
    defparam add_283_1.INJECT1_1 = "NO";
    CCU2D add_281_7 (.A0(n1025[4]), .B0(n1025[5]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n40430), 
          .S0(n1038[5]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_281_7.INIT0 = 16'h5999;
    defparam add_281_7.INIT1 = 16'h0000;
    defparam add_281_7.INJECT1_0 = "NO";
    defparam add_281_7.INJECT1_1 = "NO";
    PFUMX i38465 (.BLUT(n46334), .ALUT(n46335), .C0(akku_o_c_3), .Z(n46336));
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_299 (.A(n46051), .B(n46111), .C(n4382[1]), 
         .D(n45896), .Z(n23044)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (C))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_299.init = 16'h0f87;
    PFUMX i38309 (.BLUT(n45490), .ALUT(n45489), .C0(n45774), .Z(n45491));
    PFUMX i38463 (.BLUT(n46331), .ALUT(n46332), .C0(oprand[4]), .Z(n122_adj_511));
    LUT4 i4544_2_lut_rep_763_3_lut_4_lut_4_lut (.A(n46051), .B(n46111), 
         .C(n45_adj_356), .D(n45900), .Z(n45884)) /* synthesis lut_function=(!(A (B (C+!(D))))) */ ;
    defparam i4544_2_lut_rep_763_3_lut_4_lut_4_lut.init = 16'h7f77;
    LUT4 i31479_2_lut_3_lut_4_lut (.A(n46055), .B(n46090), .C(n6_adj_369), 
         .D(n4_adj_403), .Z(n38213)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C (D)))+!A !(C (D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i31479_2_lut_3_lut_4_lut.init = 16'h7080;
    LUT4 i2661_4_lut_4_lut (.A(n45860), .B(n45866), .C(n45864), .D(n22894), 
         .Z(n8_adj_433)) /* synthesis lut_function=(A (B+!(D))+!A !(B (D)+!B ((D)+!C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2661_4_lut_4_lut.init = 16'h88fe;
    PFUMX i38461 (.BLUT(n43557), .ALUT(n46329), .C0(akku_o_c_1), .Z(n46330));
    LUT4 mux_22_i7_3_lut_4_lut (.A(oprand[0]), .B(akku_o_c_0), .C(n16[7]), 
         .D(n16[6]), .Z(n93)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_22_i7_3_lut_4_lut.init = 16'hfe10;
    FD1P3AX oprand_i0_i2_rep_1175 (.D(data[2]), .SP(clk_c_enable_26), .CK(clk_c), 
            .Q(n46876)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam oprand_i0_i2_rep_1175.GSR = "ENABLED";
    LUT4 i31477_2_lut_3_lut_4_lut (.A(n46055), .B(n46090), .C(n6_adj_369), 
         .D(n4_adj_403), .Z(n1530[3])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(44[4] 46[11])
    defparam i31477_2_lut_3_lut_4_lut.init = 16'h8778;
    LUT4 i23869_2_lut_3_lut_4_lut (.A(n46882), .B(n46880), .C(n1156[2]), 
         .D(n43341), .Z(n545[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i23869_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i2_3_lut_4_lut_adj_300 (.A(n46882), .B(n46880), .C(akku_o_c_1), 
         .D(n46878), .Z(n23565)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut_adj_300.init = 16'hfffe;
    LUT4 i37021_2_lut_rep_997_2_lut_3_lut_4_lut (.A(n46882), .B(n46880), 
         .C(n29_adj_353), .D(n46127), .Z(n46118)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;
    defparam i37021_2_lut_rep_997_2_lut_3_lut_4_lut.init = 16'hf0f1;
    PFUMX i38457 (.BLUT(n46322), .ALUT(n46323), .C0(oprand[1]), .Z(n46324));
    LUT4 i1_2_lut_rep_1007_3_lut (.A(n46882), .B(n46880), .C(n43341), 
         .Z(n46128)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_1007_3_lut.init = 16'hfefe;
    LUT4 mux_22_i3_3_lut_4_lut (.A(n46882), .B(n46880), .C(n16[3]), .D(n16[2]), 
         .Z(n217)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_22_i3_3_lut_4_lut.init = 16'hfe10;
    PFUMX i38455 (.BLUT(n46319), .ALUT(n46320), .C0(akku_o_c_0), .Z(n122_adj_437));
    LUT4 i2254_2_lut_rep_906_3_lut_4_lut (.A(n46085), .B(n46056), .C(n4_adj_317), 
         .D(n23063), .Z(n46027)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i2254_2_lut_rep_906_3_lut_4_lut.init = 16'hffbf;
    PFUMX i38452 (.BLUT(n46315), .ALUT(n46316), .C0(oprand[0]), .Z(n122_adj_510));
    PFUMX i38177 (.BLUT(n895[0]), .ALUT(n45247), .C0(n43563), .Z(n45248));
    LUT4 mux_22_i2_3_lut_4_lut (.A(oprand[0]), .B(akku_o_c_0), .C(n16[2]), 
         .D(n16[1]), .Z(n248)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_22_i2_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_22_i1_3_lut_4_lut (.A(oprand[0]), .B(akku_o_c_0), .C(n16[1]), 
         .D(n16[0]), .Z(n159)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_22_i1_3_lut_4_lut.init = 16'hfe10;
    LUT4 i31998_2_lut_3_lut_4_lut (.A(n46057), .B(n46155), .C(n46058), 
         .D(n23881), .Z(n201[6])) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C)+!B !(C (D)+!C !(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam i31998_2_lut_3_lut_4_lut.init = 16'hb40f;
    CCU2D add_281_5 (.A0(n1025[2]), .B0(n1025[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1025[3]), .B1(n1025[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40429), .COUT(n40430), .S0(n1038[3]), .S1(n1038[4]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_281_5.INIT0 = 16'h5999;
    defparam add_281_5.INIT1 = 16'h5666;
    defparam add_281_5.INJECT1_0 = "NO";
    defparam add_281_5.INJECT1_1 = "NO";
    CCU2D add_281_3 (.A0(n1025[0]), .B0(n1025[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n1025[1]), .B1(n1025[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n40428), .COUT(n40429), .S0(n1038[1]), .S1(n1038[2]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_281_3.INIT0 = 16'h5999;
    defparam add_281_3.INIT1 = 16'h5999;
    defparam add_281_3.INJECT1_0 = "NO";
    defparam add_281_3.INJECT1_1 = "NO";
    CCU2D add_281_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n46229), .B1(n46230), .C1(n462[2]), .D1(n45904), .COUT(n40428), 
          .S1(n1038[0]));   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(45[25:40])
    defparam add_281_1.INIT0 = 16'hF000;
    defparam add_281_1.INIT1 = 16'h0e1f;
    defparam add_281_1.INJECT1_0 = "NO";
    defparam add_281_1.INJECT1_1 = "NO";
    PFUMX i38304 (.BLUT(n45479), .ALUT(n45478), .C0(oprand[3]), .Z(n45480));
    LUT4 i15820_4_lut (.A(akku_o_c_5), .B(akku_o_8__N_67[5]), .C(n46276), 
         .D(data[5]), .Z(n22547)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(73[13] 82[22])
    defparam i15820_4_lut.init = 16'hc0c5;
    FD1P3AX oprand_i0_i3_rep_1174 (.D(data[3]), .SP(clk_c_enable_26), .CK(clk_c), 
            .Q(n46875)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam oprand_i0_i3_rep_1174.GSR = "ENABLED";
    LUT4 i23836_2_lut_rep_1011_3_lut (.A(oprand[0]), .B(n46880), .C(n16[8]), 
         .Z(n46132)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i23836_2_lut_rep_1011_3_lut.init = 16'he0e0;
    FD1P3AX oprand_i0_i4_rep_1172 (.D(data[4]), .SP(clk_c_enable_26), .CK(clk_c), 
            .Q(n46873)) /* synthesis LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=18, LSE_LLINE=43, LSE_RLINE=43 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/tb02cpu2.vhd(56[9] 108[16])
    defparam oprand_i0_i4_rep_1172.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \sram64kx8("sram64kx8.dat")(1,13) 
//

module \sram64kx8("sram64kx8.dat")(1,13)  (data, address, data_7__N_89, 
            akku_o_c_4, n46211, data_7__N_102, n46237, n23757, akku_o_c_0, 
            akku_o_c_7, akku_o_c_6, akku_o_c_5, akku_o_c_3, akku_o_c_2, 
            akku_o_c_1, reset_c, clk_c, \states[0] , \states[1] );
    output [7:0]data;
    input [5:0]address;
    output [7:0]data_7__N_89;
    input akku_o_c_4;
    input n46211;
    output data_7__N_102;
    input n46237;
    input n23757;
    input akku_o_c_0;
    input akku_o_c_7;
    input akku_o_c_6;
    input akku_o_c_5;
    input akku_o_c_3;
    input akku_o_c_2;
    input akku_o_c_1;
    input reset_c;
    input clk_c;
    input \states[0] ;
    input \states[1] ;
    
    wire mem_63__7__N_297 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_63__7__N_297 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_62__7__N_294 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_62__7__N_294 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_61__7__N_291 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_61__7__N_291 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_60__7__N_288 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_60__7__N_288 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_59__7__N_285 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_59__7__N_285 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_58__7__N_282 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_58__7__N_282 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_57__7__N_279 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_57__7__N_279 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_56__7__N_276 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_56__7__N_276 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_55__7__N_273 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_55__7__N_273 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_54__7__N_270 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_54__7__N_270 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_53__7__N_267 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_53__7__N_267 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_52__7__N_264 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_52__7__N_264 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_51__7__N_261 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_51__7__N_261 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_50__7__N_258 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_50__7__N_258 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_49__7__N_255 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_49__7__N_255 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_48__7__N_252 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_48__7__N_252 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_47__7__N_249 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_47__7__N_249 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_46__7__N_246 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_46__7__N_246 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_45__7__N_243 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_45__7__N_243 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_44__7__N_240 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_44__7__N_240 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_43__7__N_237 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_43__7__N_237 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_42__7__N_234 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_42__7__N_234 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_41__7__N_231 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_41__7__N_231 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_40__7__N_228 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_40__7__N_228 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_39__7__N_225 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_39__7__N_225 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_38__7__N_222 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_38__7__N_222 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_37__7__N_219 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_37__7__N_219 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_36__7__N_216 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_36__7__N_216 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_35__7__N_213 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_35__7__N_213 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_34__7__N_210 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_34__7__N_210 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_33__7__N_207 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_33__7__N_207 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_32__7__N_204 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_32__7__N_204 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_31__7__N_201 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_31__7__N_201 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_30__7__N_198 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_30__7__N_198 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_29__7__N_195 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_29__7__N_195 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_28__7__N_192 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_28__7__N_192 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_27__7__N_189 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_27__7__N_189 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_26__7__N_186 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_26__7__N_186 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_25__7__N_183 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_25__7__N_183 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_24__7__N_180 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_24__7__N_180 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_23__7__N_177 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_23__7__N_177 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_22__7__N_174 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_22__7__N_174 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_21__7__N_171 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_21__7__N_171 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_20__7__N_168 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_20__7__N_168 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_19__7__N_165 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_19__7__N_165 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_18__7__N_162 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_18__7__N_162 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_17__7__N_159 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_17__7__N_159 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_16__7__N_156 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_16__7__N_156 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_15__7__N_153 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_15__7__N_153 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_14__7__N_150 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_14__7__N_150 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_13__7__N_147 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_13__7__N_147 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_12__7__N_144 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_12__7__N_144 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_11__7__N_141 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_11__7__N_141 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_10__7__N_138 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_10__7__N_138 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_9__7__N_135 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_9__7__N_135 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_8__7__N_132 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_8__7__N_132 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_7__7__N_129 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_7__7__N_129 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_6__7__N_126 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_6__7__N_126 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_5__7__N_123 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_5__7__N_123 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_4__7__N_120 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_4__7__N_120 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_3__7__N_117 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_3__7__N_117 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_2__7__N_114 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_2__7__N_114 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_1__7__N_111 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_1__7__N_111 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire mem_0__7__N_106 /* synthesis is_clock=1, SET_AS_NETWORK=\RAM/mem_0__7__N_106 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/cpu2system.vhd(8[13:16])
    wire [7:0]\mem[63] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[62] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[61] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[60] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[59] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[58] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[57] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[56] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[55] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[54] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[53] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[52] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[51] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[50] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[49] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[48] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[47] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[46] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[45] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[44] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[43] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[42] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[41] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[40] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[39] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[38] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[37] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[36] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[35] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[34] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[33] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[32] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[31] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[30] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[29] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[28] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[27] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[26] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[25] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[24] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[23] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[22] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[21] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[20] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[19] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[18] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[17] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[16] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[15] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[14] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[13] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[12] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[11] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[10] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[9] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[8] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[7] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[6] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[5] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[4] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[3] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[2] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[1] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    wire [7:0]\mem[0] ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(27[9:12])
    
    wire n44436, n44467, n44405, n44498, n44374, n44529, n44343, 
        n44560, n44312, n44591, n44281, n44622, n44250, n44653, 
        n44219, n44684, n44616, n44617, n44620, n44618, n44619, 
        n44621, n44647, n44648, n44651, n44649, n44650, n44652, 
        n44678, n44679, n44682, n44680, n44681, n44683, n44213, 
        n44214, n44217, n44215, n44216, n44218, n44244, n44245, 
        n44248, n44246, n44247, n44249, n44275, n44276, n44279, 
        n44277, n44278, n44280, n44492, n44493, n44496, n44494, 
        n44495, n44497, n44306, n44307, n44310, n44308, n44309, 
        n44311, n44523, n44524, n44527, n44525, n44526, n44528, 
        n44337, n44338, n44341, n44339, n44340, n44342, n44554, 
        n44555, n44558, n44556, n44557, n44559, n44368, n44369, 
        n44372, n44370, n44371, n44373, n44399, n44400, n44403, 
        n44401, n44402, n44404, n44585, n44586, n44589, n44587, 
        n44588, n44590, n44430, n44431, n44434, n44432, n44433, 
        n44435, n44461, n44462, n44465, n44463, n44464, n44466, 
        n44608, n44609, n44610, n44611, n44612, n44613, n44614, 
        n44615, n44447, n44448, n44458, n44205, n44206, n44639, 
        n44640, n44207, n44208, n44641, n44642, n44643, n44644, 
        n44645, n44646, n44209, n44210, n44670, n44671, n44672, 
        n44673, n44674, n44675, n44676, n44677, n44211, n44212, 
        n44236, n44237, n44238, n44239, n44240, n44241, n44242, 
        n44243, n44484, n44485, n44486, n44487, n44267, n44268, 
        n44269, n44270, n44271, n44272, n44273, n44274, n44488, 
        n44489, n44490, n44491, n44298, n44299, n44300, n44301, 
        n44302, n44303, n44304, n44305, n44515, n44516, n44517, 
        n44518, n44519, n44520, n44521, n44522, n44329, n44330, 
        n44331, n44332, n44333, n44334, n44335, n44336, n44546, 
        n44547, n44548, n44549, n44550, n44551, n44552, n44553, 
        n44360, n44361, n44362, n44363, n44364, n44365, n44366, 
        n44367, n44391, n44392, n44393, n44394, n44395, n44396, 
        n44397, n44398, n44577, n44578, n44579, n44580, n44581, 
        n44582, n44422, n44423, n44583, n44584, n44424, n44425, 
        n44426, n44427, n44428, n44429, n44453, n44454, n44455, 
        n44456, n44457, n44459, n44460, n44189, n44190, n46273, 
        n46236, n46238, n44191, n44192, n44449, n44450, n44193, 
        n44194, n44195, n44196, n44197, n44198, n44199, n44200, 
        n44623, n44624, n44201, n44202, n44625, n44626, n44203, 
        n44204, n44627, n44628, n46274, n44629, n44630, n46232, 
        n44631, n44632, n44633, n44634, n44635, n44636, n44637, 
        n44638, n44654, n44655, n44656, n44657, n44658, n44659, 
        n44660, n44661, n44662, n44663, n44664, n44665, n44666, 
        n44667, n44668, n44669, n44607, n44220, n44221, n44222, 
        n44223, n44224, n44225, n44226, n44227, n44228, n44229, 
        n44230, n44231, n44232, n44233, n44234, n44235, n44468, 
        n44469, n44606, n44451, n44452, n44470, n44471, n44472, 
        n44473, n44474, n44475, n44444, n44443, n44442, n44441, 
        n44440, n44439, n44251, n44252, n46239, n44605, n44604, 
        n44253, n44254, n44438, n44437, n44421, n44603, n44602, 
        n46275, n44255, n44256, n44420, n44419, n44418, n44417, 
        n44416, n44415, n44414, n44476, n44477, n44413, n44601, 
        n44412, n44600, n44576, n44575, n44411, n44410, n44409, 
        n44408, n44478, n44479, n44407, n44406, n44574, n44480, 
        n44481, n44573, n44572, n44482, n44483, n44571, n44570, 
        n44569, n44568, n44567, n44566, n44565, n44257, n44258, 
        n44564, n44563, n44562, n44561, n44390, n44389, n44388, 
        n44387, n44386, n44385, n44384, n44383, n44259, n44260, 
        n44261, n44262, n44382, n44263, n44264, n44381, n44592, 
        n44593, n44380, n44379, n44378, n44265, n44266, n44377, 
        n44376, n44375, n44359, n44358, n44357, n44499, n44500, 
        n44356, n44355, n44354, n44353, n44352, n44351, n44350, 
        n44349, n44348, n44347, n44346, n44282, n44283, n44345, 
        n44344, n44545, n44544, n44284, n44285, n44501, n44502, 
        n44543, n44542, n44541, n44286, n44287, n44599, n44540, 
        n44539, n44538, n44537, n44536, n44598, n44535, n44534, 
        n44533, n44532, n44531, n44530, n44328, n44327, n44326, 
        n44325, n44288, n44289, n44324, n44323, n44290, n44291, 
        n44322, n44321, n44320, n44597, n44319, n44292, n44293, 
        n44594, n44595, n44294, n44295, n44318, n44317, n44296, 
        n44297, n44503, n44504, n46234, n44316, n44315, n44596, 
        n44314, n44505, n44506, n44313, n44514, n44513, n44512, 
        n44511, n44507, n44508, n44510, n46241, n44509, n44445, 
        n44446, n46856, n43653, n46220, n43635, n46242, n43636, 
        n43654, n46172, n46278;
    
    FD1S1A data_7__I_0_i1 (.D(data[0]), .CK(mem_63__7__N_297), .Q(\mem[63] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5187_i1 (.D(data[0]), .CK(mem_62__7__N_294), .Q(\mem[62] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i1 (.D(data[0]), .CK(mem_61__7__N_291), .Q(\mem[61] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i1 (.D(data[0]), .CK(mem_60__7__N_288), .Q(\mem[60] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i1 (.D(data[0]), .CK(mem_59__7__N_285), .Q(\mem[59] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i1 (.D(data[0]), .CK(mem_58__7__N_282), .Q(\mem[58] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i1 (.D(data[0]), .CK(mem_57__7__N_279), .Q(\mem[57] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i1 (.D(data[0]), .CK(mem_56__7__N_276), .Q(\mem[56] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i1 (.D(data[0]), .CK(mem_55__7__N_273), .Q(\mem[55] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i1 (.D(data[0]), .CK(mem_54__7__N_270), .Q(\mem[54] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i1 (.D(data[0]), .CK(mem_53__7__N_267), .Q(\mem[53] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i1 (.D(data[0]), .CK(mem_52__7__N_264), .Q(\mem[52] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i1 (.D(data[0]), .CK(mem_51__7__N_261), .Q(\mem[51] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i1 (.D(data[0]), .CK(mem_50__7__N_258), .Q(\mem[50] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i1 (.D(data[0]), .CK(mem_49__7__N_255), .Q(\mem[49] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i1 (.D(data[0]), .CK(mem_48__7__N_252), .Q(\mem[48] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i1 (.D(data[0]), .CK(mem_47__7__N_249), .Q(\mem[47] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i1 (.D(data[0]), .CK(mem_46__7__N_246), .Q(\mem[46] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i1 (.D(data[0]), .CK(mem_45__7__N_243), .Q(\mem[45] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i1 (.D(data[0]), .CK(mem_44__7__N_240), .Q(\mem[44] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i1 (.D(data[0]), .CK(mem_43__7__N_237), .Q(\mem[43] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i1 (.D(data[0]), .CK(mem_42__7__N_234), .Q(\mem[42] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i1 (.D(data[0]), .CK(mem_41__7__N_231), .Q(\mem[41] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i1 (.D(data[0]), .CK(mem_40__7__N_228), .Q(\mem[40] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i1 (.D(data[0]), .CK(mem_39__7__N_225), .Q(\mem[39] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i1 (.D(data[0]), .CK(mem_38__7__N_222), .Q(\mem[38] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i1 (.D(data[0]), .CK(mem_37__7__N_219), .Q(\mem[37] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i1 (.D(data[0]), .CK(mem_36__7__N_216), .Q(\mem[36] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i1 (.D(data[0]), .CK(mem_35__7__N_213), .Q(\mem[35] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i1 (.D(data[0]), .CK(mem_34__7__N_210), .Q(\mem[34] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i1 (.D(data[0]), .CK(mem_33__7__N_207), .Q(\mem[33] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i1 (.D(data[0]), .CK(mem_32__7__N_204), .Q(\mem[32] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i1 (.D(data[0]), .CK(mem_31__7__N_201), .Q(\mem[31] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i1 (.D(data[0]), .CK(mem_30__7__N_198), .Q(\mem[30] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i1 (.D(data[0]), .CK(mem_29__7__N_195), .Q(\mem[29] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i1 (.D(data[0]), .CK(mem_28__7__N_192), .Q(\mem[28] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i1 (.D(data[0]), .CK(mem_27__7__N_189), .Q(\mem[27] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i1 (.D(data[0]), .CK(mem_26__7__N_186), .Q(\mem[26] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i1 (.D(data[0]), .CK(mem_25__7__N_183), .Q(\mem[25] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i1 (.D(data[0]), .CK(mem_24__7__N_180), .Q(\mem[24] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i1 (.D(data[0]), .CK(mem_23__7__N_177), .Q(\mem[23] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i1 (.D(data[0]), .CK(mem_22__7__N_174), .Q(\mem[22] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i1 (.D(data[0]), .CK(mem_21__7__N_171), .Q(\mem[21] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5061_i1 (.D(data[0]), .CK(mem_20__7__N_168), .Q(\mem[20] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i1 (.D(data[0]), .CK(mem_19__7__N_165), .Q(\mem[19] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5055_i1 (.D(data[0]), .CK(mem_18__7__N_162), .Q(\mem[18] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5052_i1 (.D(data[0]), .CK(mem_17__7__N_159), .Q(\mem[17] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i1 (.D(data[0]), .CK(mem_16__7__N_156), .Q(\mem[16] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5046_i1 (.D(data[0]), .CK(mem_15__7__N_153), .Q(\mem[15] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5043_i1 (.D(data[0]), .CK(mem_14__7__N_150), .Q(\mem[14] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5040_i1 (.D(data[0]), .CK(mem_13__7__N_147), .Q(\mem[13] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5037_i1 (.D(data[0]), .CK(mem_12__7__N_144), .Q(\mem[12] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i1 (.D(data[0]), .CK(mem_11__7__N_141), .Q(\mem[11] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5031_i1 (.D(data[0]), .CK(mem_10__7__N_138), .Q(\mem[10] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5028_i1 (.D(data[0]), .CK(mem_9__7__N_135), .Q(\mem[9] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5025_i1 (.D(data[0]), .CK(mem_8__7__N_132), .Q(\mem[8] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5022_i1 (.D(data[0]), .CK(mem_7__7__N_129), .Q(\mem[7] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5019_i1 (.D(data[0]), .CK(mem_6__7__N_126), .Q(\mem[6] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5016_i1 (.D(data[0]), .CK(mem_5__7__N_123), .Q(\mem[5] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5013_i1 (.D(data[0]), .CK(mem_4__7__N_120), .Q(\mem[4] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5010_i1 (.D(data[0]), .CK(mem_3__7__N_117), .Q(\mem[3] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i1.GSR = "DISABLED";
    FD1S1A data_7__I_0_5007_i1 (.D(data[0]), .CK(mem_2__7__N_114), .Q(\mem[2] [0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i1.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5004_i1 (.D(data[0]), .CK(mem_1__7__N_111), .Q(\mem[1] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i1.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5002_i1 (.D(data[0]), .CK(mem_0__7__N_106), .Q(\mem[0] [0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i1.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5002_i2 (.D(data[1]), .CK(mem_0__7__N_106), .Q(\mem[0] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5002_i3 (.D(data[2]), .CK(mem_0__7__N_106), .Q(\mem[0] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5002_i4 (.D(data[3]), .CK(mem_0__7__N_106), .Q(\mem[0] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5002_i5 (.D(data[4]), .CK(mem_0__7__N_106), .Q(\mem[0] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i5.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5002_i6 (.D(data[5]), .CK(mem_0__7__N_106), .Q(\mem[0] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5002_i7 (.D(data[6]), .CK(mem_0__7__N_106), .Q(\mem[0] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i7.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5002_i8 (.D(data[7]), .CK(mem_0__7__N_106), .Q(\mem[0] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5002_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5004_i2 (.D(data[1]), .CK(mem_1__7__N_111), .Q(\mem[1] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i2.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5004_i3 (.D(data[2]), .CK(mem_1__7__N_111), .Q(\mem[1] [2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5004_i4 (.D(data[3]), .CK(mem_1__7__N_111), .Q(\mem[1] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5004_i5 (.D(data[4]), .CK(mem_1__7__N_111), .Q(\mem[1] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i5.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5004_i6 (.D(data[5]), .CK(mem_1__7__N_111), .Q(\mem[1] [5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i6.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5004_i7 (.D(data[6]), .CK(mem_1__7__N_111), .Q(\mem[1] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i7.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5004_i8 (.D(data[7]), .CK(mem_1__7__N_111), .Q(\mem[1] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5004_i8.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5007_i2 (.D(data[1]), .CK(mem_2__7__N_114), .Q(\mem[2] [1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5007_i3 (.D(data[2]), .CK(mem_2__7__N_114), .Q(\mem[2] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5007_i4 (.D(data[3]), .CK(mem_2__7__N_114), .Q(\mem[2] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5007_i5 (.D(data[4]), .CK(mem_2__7__N_114), .Q(\mem[2] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5007_i6 (.D(data[5]), .CK(mem_2__7__N_114), .Q(\mem[2] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i6.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5007_i7 (.D(data[6]), .CK(mem_2__7__N_114), .Q(\mem[2] [6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i7.GSR = "DISABLED";
    FD1S1AY data_7__I_0_5007_i8 (.D(data[7]), .CK(mem_2__7__N_114), .Q(\mem[2] [7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5007_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_i2 (.D(data[1]), .CK(mem_63__7__N_297), .Q(\mem[63] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_i3 (.D(data[2]), .CK(mem_63__7__N_297), .Q(\mem[63] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_i4 (.D(data[3]), .CK(mem_63__7__N_297), .Q(\mem[63] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_i5 (.D(data[4]), .CK(mem_63__7__N_297), .Q(\mem[63] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_i6 (.D(data[5]), .CK(mem_63__7__N_297), .Q(\mem[63] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_i7 (.D(data[6]), .CK(mem_63__7__N_297), .Q(\mem[63] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_i8 (.D(data[7]), .CK(mem_63__7__N_297), .Q(\mem[63] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5187_i2 (.D(data[1]), .CK(mem_62__7__N_294), .Q(\mem[62] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5187_i3 (.D(data[2]), .CK(mem_62__7__N_294), .Q(\mem[62] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5187_i4 (.D(data[3]), .CK(mem_62__7__N_294), .Q(\mem[62] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5187_i5 (.D(data[4]), .CK(mem_62__7__N_294), .Q(\mem[62] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5187_i6 (.D(data[5]), .CK(mem_62__7__N_294), .Q(\mem[62] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5187_i7 (.D(data[6]), .CK(mem_62__7__N_294), .Q(\mem[62] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5187_i8 (.D(data[7]), .CK(mem_62__7__N_294), .Q(\mem[62] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5187_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i2 (.D(data[1]), .CK(mem_61__7__N_291), .Q(\mem[61] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i3 (.D(data[2]), .CK(mem_61__7__N_291), .Q(\mem[61] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i4 (.D(data[3]), .CK(mem_61__7__N_291), .Q(\mem[61] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i5 (.D(data[4]), .CK(mem_61__7__N_291), .Q(\mem[61] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i6 (.D(data[5]), .CK(mem_61__7__N_291), .Q(\mem[61] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i7 (.D(data[6]), .CK(mem_61__7__N_291), .Q(\mem[61] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5184_i8 (.D(data[7]), .CK(mem_61__7__N_291), .Q(\mem[61] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5184_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i2 (.D(data[1]), .CK(mem_60__7__N_288), .Q(\mem[60] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i3 (.D(data[2]), .CK(mem_60__7__N_288), .Q(\mem[60] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i4 (.D(data[3]), .CK(mem_60__7__N_288), .Q(\mem[60] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i5 (.D(data[4]), .CK(mem_60__7__N_288), .Q(\mem[60] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i6 (.D(data[5]), .CK(mem_60__7__N_288), .Q(\mem[60] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i7 (.D(data[6]), .CK(mem_60__7__N_288), .Q(\mem[60] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5181_i8 (.D(data[7]), .CK(mem_60__7__N_288), .Q(\mem[60] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5181_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i2 (.D(data[1]), .CK(mem_59__7__N_285), .Q(\mem[59] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i3 (.D(data[2]), .CK(mem_59__7__N_285), .Q(\mem[59] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i4 (.D(data[3]), .CK(mem_59__7__N_285), .Q(\mem[59] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i5 (.D(data[4]), .CK(mem_59__7__N_285), .Q(\mem[59] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i6 (.D(data[5]), .CK(mem_59__7__N_285), .Q(\mem[59] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i7 (.D(data[6]), .CK(mem_59__7__N_285), .Q(\mem[59] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5178_i8 (.D(data[7]), .CK(mem_59__7__N_285), .Q(\mem[59] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5178_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i2 (.D(data[1]), .CK(mem_58__7__N_282), .Q(\mem[58] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i3 (.D(data[2]), .CK(mem_58__7__N_282), .Q(\mem[58] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i4 (.D(data[3]), .CK(mem_58__7__N_282), .Q(\mem[58] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i5 (.D(data[4]), .CK(mem_58__7__N_282), .Q(\mem[58] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i6 (.D(data[5]), .CK(mem_58__7__N_282), .Q(\mem[58] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i7 (.D(data[6]), .CK(mem_58__7__N_282), .Q(\mem[58] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5175_i8 (.D(data[7]), .CK(mem_58__7__N_282), .Q(\mem[58] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5175_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i2 (.D(data[1]), .CK(mem_57__7__N_279), .Q(\mem[57] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i3 (.D(data[2]), .CK(mem_57__7__N_279), .Q(\mem[57] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i4 (.D(data[3]), .CK(mem_57__7__N_279), .Q(\mem[57] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i5 (.D(data[4]), .CK(mem_57__7__N_279), .Q(\mem[57] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i6 (.D(data[5]), .CK(mem_57__7__N_279), .Q(\mem[57] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i7 (.D(data[6]), .CK(mem_57__7__N_279), .Q(\mem[57] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5172_i8 (.D(data[7]), .CK(mem_57__7__N_279), .Q(\mem[57] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5172_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i2 (.D(data[1]), .CK(mem_56__7__N_276), .Q(\mem[56] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i3 (.D(data[2]), .CK(mem_56__7__N_276), .Q(\mem[56] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i4 (.D(data[3]), .CK(mem_56__7__N_276), .Q(\mem[56] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i5 (.D(data[4]), .CK(mem_56__7__N_276), .Q(\mem[56] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i6 (.D(data[5]), .CK(mem_56__7__N_276), .Q(\mem[56] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i7 (.D(data[6]), .CK(mem_56__7__N_276), .Q(\mem[56] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5169_i8 (.D(data[7]), .CK(mem_56__7__N_276), .Q(\mem[56] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5169_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i2 (.D(data[1]), .CK(mem_55__7__N_273), .Q(\mem[55] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i3 (.D(data[2]), .CK(mem_55__7__N_273), .Q(\mem[55] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i4 (.D(data[3]), .CK(mem_55__7__N_273), .Q(\mem[55] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i5 (.D(data[4]), .CK(mem_55__7__N_273), .Q(\mem[55] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i6 (.D(data[5]), .CK(mem_55__7__N_273), .Q(\mem[55] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i7 (.D(data[6]), .CK(mem_55__7__N_273), .Q(\mem[55] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5166_i8 (.D(data[7]), .CK(mem_55__7__N_273), .Q(\mem[55] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5166_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i2 (.D(data[1]), .CK(mem_54__7__N_270), .Q(\mem[54] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i3 (.D(data[2]), .CK(mem_54__7__N_270), .Q(\mem[54] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i4 (.D(data[3]), .CK(mem_54__7__N_270), .Q(\mem[54] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i5 (.D(data[4]), .CK(mem_54__7__N_270), .Q(\mem[54] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i6 (.D(data[5]), .CK(mem_54__7__N_270), .Q(\mem[54] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i7 (.D(data[6]), .CK(mem_54__7__N_270), .Q(\mem[54] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5163_i8 (.D(data[7]), .CK(mem_54__7__N_270), .Q(\mem[54] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5163_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i2 (.D(data[1]), .CK(mem_53__7__N_267), .Q(\mem[53] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i3 (.D(data[2]), .CK(mem_53__7__N_267), .Q(\mem[53] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i4 (.D(data[3]), .CK(mem_53__7__N_267), .Q(\mem[53] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i5 (.D(data[4]), .CK(mem_53__7__N_267), .Q(\mem[53] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i6 (.D(data[5]), .CK(mem_53__7__N_267), .Q(\mem[53] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i7 (.D(data[6]), .CK(mem_53__7__N_267), .Q(\mem[53] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5160_i8 (.D(data[7]), .CK(mem_53__7__N_267), .Q(\mem[53] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5160_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i2 (.D(data[1]), .CK(mem_52__7__N_264), .Q(\mem[52] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i3 (.D(data[2]), .CK(mem_52__7__N_264), .Q(\mem[52] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i4 (.D(data[3]), .CK(mem_52__7__N_264), .Q(\mem[52] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i5 (.D(data[4]), .CK(mem_52__7__N_264), .Q(\mem[52] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i6 (.D(data[5]), .CK(mem_52__7__N_264), .Q(\mem[52] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i7 (.D(data[6]), .CK(mem_52__7__N_264), .Q(\mem[52] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5157_i8 (.D(data[7]), .CK(mem_52__7__N_264), .Q(\mem[52] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5157_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i2 (.D(data[1]), .CK(mem_51__7__N_261), .Q(\mem[51] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i3 (.D(data[2]), .CK(mem_51__7__N_261), .Q(\mem[51] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i4 (.D(data[3]), .CK(mem_51__7__N_261), .Q(\mem[51] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i5 (.D(data[4]), .CK(mem_51__7__N_261), .Q(\mem[51] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i6 (.D(data[5]), .CK(mem_51__7__N_261), .Q(\mem[51] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i7 (.D(data[6]), .CK(mem_51__7__N_261), .Q(\mem[51] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5154_i8 (.D(data[7]), .CK(mem_51__7__N_261), .Q(\mem[51] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5154_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i2 (.D(data[1]), .CK(mem_50__7__N_258), .Q(\mem[50] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i3 (.D(data[2]), .CK(mem_50__7__N_258), .Q(\mem[50] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i4 (.D(data[3]), .CK(mem_50__7__N_258), .Q(\mem[50] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i5 (.D(data[4]), .CK(mem_50__7__N_258), .Q(\mem[50] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i6 (.D(data[5]), .CK(mem_50__7__N_258), .Q(\mem[50] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i7 (.D(data[6]), .CK(mem_50__7__N_258), .Q(\mem[50] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5151_i8 (.D(data[7]), .CK(mem_50__7__N_258), .Q(\mem[50] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5151_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i2 (.D(data[1]), .CK(mem_49__7__N_255), .Q(\mem[49] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i3 (.D(data[2]), .CK(mem_49__7__N_255), .Q(\mem[49] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i4 (.D(data[3]), .CK(mem_49__7__N_255), .Q(\mem[49] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i5 (.D(data[4]), .CK(mem_49__7__N_255), .Q(\mem[49] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i6 (.D(data[5]), .CK(mem_49__7__N_255), .Q(\mem[49] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i7 (.D(data[6]), .CK(mem_49__7__N_255), .Q(\mem[49] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5148_i8 (.D(data[7]), .CK(mem_49__7__N_255), .Q(\mem[49] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5148_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i2 (.D(data[1]), .CK(mem_48__7__N_252), .Q(\mem[48] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i3 (.D(data[2]), .CK(mem_48__7__N_252), .Q(\mem[48] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i4 (.D(data[3]), .CK(mem_48__7__N_252), .Q(\mem[48] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i5 (.D(data[4]), .CK(mem_48__7__N_252), .Q(\mem[48] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i6 (.D(data[5]), .CK(mem_48__7__N_252), .Q(\mem[48] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i7 (.D(data[6]), .CK(mem_48__7__N_252), .Q(\mem[48] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5145_i8 (.D(data[7]), .CK(mem_48__7__N_252), .Q(\mem[48] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5145_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i2 (.D(data[1]), .CK(mem_47__7__N_249), .Q(\mem[47] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i3 (.D(data[2]), .CK(mem_47__7__N_249), .Q(\mem[47] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i4 (.D(data[3]), .CK(mem_47__7__N_249), .Q(\mem[47] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i5 (.D(data[4]), .CK(mem_47__7__N_249), .Q(\mem[47] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i6 (.D(data[5]), .CK(mem_47__7__N_249), .Q(\mem[47] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i7 (.D(data[6]), .CK(mem_47__7__N_249), .Q(\mem[47] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5142_i8 (.D(data[7]), .CK(mem_47__7__N_249), .Q(\mem[47] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5142_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i2 (.D(data[1]), .CK(mem_46__7__N_246), .Q(\mem[46] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i3 (.D(data[2]), .CK(mem_46__7__N_246), .Q(\mem[46] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i4 (.D(data[3]), .CK(mem_46__7__N_246), .Q(\mem[46] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i5 (.D(data[4]), .CK(mem_46__7__N_246), .Q(\mem[46] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i6 (.D(data[5]), .CK(mem_46__7__N_246), .Q(\mem[46] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i7 (.D(data[6]), .CK(mem_46__7__N_246), .Q(\mem[46] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5139_i8 (.D(data[7]), .CK(mem_46__7__N_246), .Q(\mem[46] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5139_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i2 (.D(data[1]), .CK(mem_45__7__N_243), .Q(\mem[45] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i3 (.D(data[2]), .CK(mem_45__7__N_243), .Q(\mem[45] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i4 (.D(data[3]), .CK(mem_45__7__N_243), .Q(\mem[45] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i5 (.D(data[4]), .CK(mem_45__7__N_243), .Q(\mem[45] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i6 (.D(data[5]), .CK(mem_45__7__N_243), .Q(\mem[45] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i7 (.D(data[6]), .CK(mem_45__7__N_243), .Q(\mem[45] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5136_i8 (.D(data[7]), .CK(mem_45__7__N_243), .Q(\mem[45] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5136_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i2 (.D(data[1]), .CK(mem_44__7__N_240), .Q(\mem[44] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i3 (.D(data[2]), .CK(mem_44__7__N_240), .Q(\mem[44] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i4 (.D(data[3]), .CK(mem_44__7__N_240), .Q(\mem[44] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i5 (.D(data[4]), .CK(mem_44__7__N_240), .Q(\mem[44] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i6 (.D(data[5]), .CK(mem_44__7__N_240), .Q(\mem[44] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i7 (.D(data[6]), .CK(mem_44__7__N_240), .Q(\mem[44] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5133_i8 (.D(data[7]), .CK(mem_44__7__N_240), .Q(\mem[44] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5133_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i2 (.D(data[1]), .CK(mem_43__7__N_237), .Q(\mem[43] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i3 (.D(data[2]), .CK(mem_43__7__N_237), .Q(\mem[43] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i4 (.D(data[3]), .CK(mem_43__7__N_237), .Q(\mem[43] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i5 (.D(data[4]), .CK(mem_43__7__N_237), .Q(\mem[43] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i6 (.D(data[5]), .CK(mem_43__7__N_237), .Q(\mem[43] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i7 (.D(data[6]), .CK(mem_43__7__N_237), .Q(\mem[43] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5130_i8 (.D(data[7]), .CK(mem_43__7__N_237), .Q(\mem[43] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5130_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i2 (.D(data[1]), .CK(mem_42__7__N_234), .Q(\mem[42] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i3 (.D(data[2]), .CK(mem_42__7__N_234), .Q(\mem[42] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i4 (.D(data[3]), .CK(mem_42__7__N_234), .Q(\mem[42] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i5 (.D(data[4]), .CK(mem_42__7__N_234), .Q(\mem[42] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i6 (.D(data[5]), .CK(mem_42__7__N_234), .Q(\mem[42] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i7 (.D(data[6]), .CK(mem_42__7__N_234), .Q(\mem[42] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5127_i8 (.D(data[7]), .CK(mem_42__7__N_234), .Q(\mem[42] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5127_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i2 (.D(data[1]), .CK(mem_41__7__N_231), .Q(\mem[41] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i3 (.D(data[2]), .CK(mem_41__7__N_231), .Q(\mem[41] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i4 (.D(data[3]), .CK(mem_41__7__N_231), .Q(\mem[41] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i5 (.D(data[4]), .CK(mem_41__7__N_231), .Q(\mem[41] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i6 (.D(data[5]), .CK(mem_41__7__N_231), .Q(\mem[41] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i7 (.D(data[6]), .CK(mem_41__7__N_231), .Q(\mem[41] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5124_i8 (.D(data[7]), .CK(mem_41__7__N_231), .Q(\mem[41] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5124_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i2 (.D(data[1]), .CK(mem_40__7__N_228), .Q(\mem[40] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i3 (.D(data[2]), .CK(mem_40__7__N_228), .Q(\mem[40] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i4 (.D(data[3]), .CK(mem_40__7__N_228), .Q(\mem[40] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i5 (.D(data[4]), .CK(mem_40__7__N_228), .Q(\mem[40] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i6 (.D(data[5]), .CK(mem_40__7__N_228), .Q(\mem[40] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i7 (.D(data[6]), .CK(mem_40__7__N_228), .Q(\mem[40] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5121_i8 (.D(data[7]), .CK(mem_40__7__N_228), .Q(\mem[40] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5121_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i2 (.D(data[1]), .CK(mem_39__7__N_225), .Q(\mem[39] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i3 (.D(data[2]), .CK(mem_39__7__N_225), .Q(\mem[39] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i4 (.D(data[3]), .CK(mem_39__7__N_225), .Q(\mem[39] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i5 (.D(data[4]), .CK(mem_39__7__N_225), .Q(\mem[39] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i6 (.D(data[5]), .CK(mem_39__7__N_225), .Q(\mem[39] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i7 (.D(data[6]), .CK(mem_39__7__N_225), .Q(\mem[39] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5118_i8 (.D(data[7]), .CK(mem_39__7__N_225), .Q(\mem[39] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5118_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i2 (.D(data[1]), .CK(mem_38__7__N_222), .Q(\mem[38] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i3 (.D(data[2]), .CK(mem_38__7__N_222), .Q(\mem[38] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i4 (.D(data[3]), .CK(mem_38__7__N_222), .Q(\mem[38] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i5 (.D(data[4]), .CK(mem_38__7__N_222), .Q(\mem[38] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i6 (.D(data[5]), .CK(mem_38__7__N_222), .Q(\mem[38] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i7 (.D(data[6]), .CK(mem_38__7__N_222), .Q(\mem[38] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5115_i8 (.D(data[7]), .CK(mem_38__7__N_222), .Q(\mem[38] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5115_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i2 (.D(data[1]), .CK(mem_37__7__N_219), .Q(\mem[37] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i3 (.D(data[2]), .CK(mem_37__7__N_219), .Q(\mem[37] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i4 (.D(data[3]), .CK(mem_37__7__N_219), .Q(\mem[37] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i5 (.D(data[4]), .CK(mem_37__7__N_219), .Q(\mem[37] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i6 (.D(data[5]), .CK(mem_37__7__N_219), .Q(\mem[37] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i7 (.D(data[6]), .CK(mem_37__7__N_219), .Q(\mem[37] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5112_i8 (.D(data[7]), .CK(mem_37__7__N_219), .Q(\mem[37] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5112_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i2 (.D(data[1]), .CK(mem_36__7__N_216), .Q(\mem[36] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i3 (.D(data[2]), .CK(mem_36__7__N_216), .Q(\mem[36] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i4 (.D(data[3]), .CK(mem_36__7__N_216), .Q(\mem[36] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i5 (.D(data[4]), .CK(mem_36__7__N_216), .Q(\mem[36] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i6 (.D(data[5]), .CK(mem_36__7__N_216), .Q(\mem[36] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i7 (.D(data[6]), .CK(mem_36__7__N_216), .Q(\mem[36] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5109_i8 (.D(data[7]), .CK(mem_36__7__N_216), .Q(\mem[36] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5109_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i2 (.D(data[1]), .CK(mem_35__7__N_213), .Q(\mem[35] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i3 (.D(data[2]), .CK(mem_35__7__N_213), .Q(\mem[35] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i4 (.D(data[3]), .CK(mem_35__7__N_213), .Q(\mem[35] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i5 (.D(data[4]), .CK(mem_35__7__N_213), .Q(\mem[35] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i6 (.D(data[5]), .CK(mem_35__7__N_213), .Q(\mem[35] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i7 (.D(data[6]), .CK(mem_35__7__N_213), .Q(\mem[35] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5106_i8 (.D(data[7]), .CK(mem_35__7__N_213), .Q(\mem[35] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5106_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i2 (.D(data[1]), .CK(mem_34__7__N_210), .Q(\mem[34] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i3 (.D(data[2]), .CK(mem_34__7__N_210), .Q(\mem[34] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i4 (.D(data[3]), .CK(mem_34__7__N_210), .Q(\mem[34] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i5 (.D(data[4]), .CK(mem_34__7__N_210), .Q(\mem[34] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i6 (.D(data[5]), .CK(mem_34__7__N_210), .Q(\mem[34] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i7 (.D(data[6]), .CK(mem_34__7__N_210), .Q(\mem[34] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5103_i8 (.D(data[7]), .CK(mem_34__7__N_210), .Q(\mem[34] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5103_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i2 (.D(data[1]), .CK(mem_33__7__N_207), .Q(\mem[33] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i3 (.D(data[2]), .CK(mem_33__7__N_207), .Q(\mem[33] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i4 (.D(data[3]), .CK(mem_33__7__N_207), .Q(\mem[33] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i5 (.D(data[4]), .CK(mem_33__7__N_207), .Q(\mem[33] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i6 (.D(data[5]), .CK(mem_33__7__N_207), .Q(\mem[33] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i7 (.D(data[6]), .CK(mem_33__7__N_207), .Q(\mem[33] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5100_i8 (.D(data[7]), .CK(mem_33__7__N_207), .Q(\mem[33] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5100_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i2 (.D(data[1]), .CK(mem_32__7__N_204), .Q(\mem[32] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i3 (.D(data[2]), .CK(mem_32__7__N_204), .Q(\mem[32] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i4 (.D(data[3]), .CK(mem_32__7__N_204), .Q(\mem[32] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i5 (.D(data[4]), .CK(mem_32__7__N_204), .Q(\mem[32] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i6 (.D(data[5]), .CK(mem_32__7__N_204), .Q(\mem[32] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i7 (.D(data[6]), .CK(mem_32__7__N_204), .Q(\mem[32] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5097_i8 (.D(data[7]), .CK(mem_32__7__N_204), .Q(\mem[32] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5097_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i2 (.D(data[1]), .CK(mem_31__7__N_201), .Q(\mem[31] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i3 (.D(data[2]), .CK(mem_31__7__N_201), .Q(\mem[31] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i4 (.D(data[3]), .CK(mem_31__7__N_201), .Q(\mem[31] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i5 (.D(data[4]), .CK(mem_31__7__N_201), .Q(\mem[31] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i6 (.D(data[5]), .CK(mem_31__7__N_201), .Q(\mem[31] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i7 (.D(data[6]), .CK(mem_31__7__N_201), .Q(\mem[31] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5094_i8 (.D(data[7]), .CK(mem_31__7__N_201), .Q(\mem[31] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5094_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i2 (.D(data[1]), .CK(mem_30__7__N_198), .Q(\mem[30] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i3 (.D(data[2]), .CK(mem_30__7__N_198), .Q(\mem[30] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i4 (.D(data[3]), .CK(mem_30__7__N_198), .Q(\mem[30] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i5 (.D(data[4]), .CK(mem_30__7__N_198), .Q(\mem[30] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i6 (.D(data[5]), .CK(mem_30__7__N_198), .Q(\mem[30] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i7 (.D(data[6]), .CK(mem_30__7__N_198), .Q(\mem[30] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5091_i8 (.D(data[7]), .CK(mem_30__7__N_198), .Q(\mem[30] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5091_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i2 (.D(data[1]), .CK(mem_29__7__N_195), .Q(\mem[29] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i3 (.D(data[2]), .CK(mem_29__7__N_195), .Q(\mem[29] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i4 (.D(data[3]), .CK(mem_29__7__N_195), .Q(\mem[29] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i5 (.D(data[4]), .CK(mem_29__7__N_195), .Q(\mem[29] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i6 (.D(data[5]), .CK(mem_29__7__N_195), .Q(\mem[29] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i7 (.D(data[6]), .CK(mem_29__7__N_195), .Q(\mem[29] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5088_i8 (.D(data[7]), .CK(mem_29__7__N_195), .Q(\mem[29] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5088_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i2 (.D(data[1]), .CK(mem_28__7__N_192), .Q(\mem[28] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i3 (.D(data[2]), .CK(mem_28__7__N_192), .Q(\mem[28] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i4 (.D(data[3]), .CK(mem_28__7__N_192), .Q(\mem[28] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i5 (.D(data[4]), .CK(mem_28__7__N_192), .Q(\mem[28] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i6 (.D(data[5]), .CK(mem_28__7__N_192), .Q(\mem[28] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i7 (.D(data[6]), .CK(mem_28__7__N_192), .Q(\mem[28] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5085_i8 (.D(data[7]), .CK(mem_28__7__N_192), .Q(\mem[28] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5085_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i2 (.D(data[1]), .CK(mem_27__7__N_189), .Q(\mem[27] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i3 (.D(data[2]), .CK(mem_27__7__N_189), .Q(\mem[27] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i4 (.D(data[3]), .CK(mem_27__7__N_189), .Q(\mem[27] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i5 (.D(data[4]), .CK(mem_27__7__N_189), .Q(\mem[27] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i6 (.D(data[5]), .CK(mem_27__7__N_189), .Q(\mem[27] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i7 (.D(data[6]), .CK(mem_27__7__N_189), .Q(\mem[27] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5082_i8 (.D(data[7]), .CK(mem_27__7__N_189), .Q(\mem[27] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5082_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i2 (.D(data[1]), .CK(mem_26__7__N_186), .Q(\mem[26] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i3 (.D(data[2]), .CK(mem_26__7__N_186), .Q(\mem[26] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i4 (.D(data[3]), .CK(mem_26__7__N_186), .Q(\mem[26] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i5 (.D(data[4]), .CK(mem_26__7__N_186), .Q(\mem[26] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i6 (.D(data[5]), .CK(mem_26__7__N_186), .Q(\mem[26] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i7 (.D(data[6]), .CK(mem_26__7__N_186), .Q(\mem[26] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5079_i8 (.D(data[7]), .CK(mem_26__7__N_186), .Q(\mem[26] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5079_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i2 (.D(data[1]), .CK(mem_25__7__N_183), .Q(\mem[25] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i3 (.D(data[2]), .CK(mem_25__7__N_183), .Q(\mem[25] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i4 (.D(data[3]), .CK(mem_25__7__N_183), .Q(\mem[25] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i5 (.D(data[4]), .CK(mem_25__7__N_183), .Q(\mem[25] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i6 (.D(data[5]), .CK(mem_25__7__N_183), .Q(\mem[25] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i7 (.D(data[6]), .CK(mem_25__7__N_183), .Q(\mem[25] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5076_i8 (.D(data[7]), .CK(mem_25__7__N_183), .Q(\mem[25] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5076_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i2 (.D(data[1]), .CK(mem_24__7__N_180), .Q(\mem[24] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i3 (.D(data[2]), .CK(mem_24__7__N_180), .Q(\mem[24] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i4 (.D(data[3]), .CK(mem_24__7__N_180), .Q(\mem[24] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i5 (.D(data[4]), .CK(mem_24__7__N_180), .Q(\mem[24] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i6 (.D(data[5]), .CK(mem_24__7__N_180), .Q(\mem[24] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i7 (.D(data[6]), .CK(mem_24__7__N_180), .Q(\mem[24] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5073_i8 (.D(data[7]), .CK(mem_24__7__N_180), .Q(\mem[24] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5073_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i2 (.D(data[1]), .CK(mem_23__7__N_177), .Q(\mem[23] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i3 (.D(data[2]), .CK(mem_23__7__N_177), .Q(\mem[23] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i4 (.D(data[3]), .CK(mem_23__7__N_177), .Q(\mem[23] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i5 (.D(data[4]), .CK(mem_23__7__N_177), .Q(\mem[23] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i6 (.D(data[5]), .CK(mem_23__7__N_177), .Q(\mem[23] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i7 (.D(data[6]), .CK(mem_23__7__N_177), .Q(\mem[23] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5070_i8 (.D(data[7]), .CK(mem_23__7__N_177), .Q(\mem[23] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5070_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i2 (.D(data[1]), .CK(mem_22__7__N_174), .Q(\mem[22] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i3 (.D(data[2]), .CK(mem_22__7__N_174), .Q(\mem[22] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i4 (.D(data[3]), .CK(mem_22__7__N_174), .Q(\mem[22] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i5 (.D(data[4]), .CK(mem_22__7__N_174), .Q(\mem[22] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i6 (.D(data[5]), .CK(mem_22__7__N_174), .Q(\mem[22] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i7 (.D(data[6]), .CK(mem_22__7__N_174), .Q(\mem[22] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5067_i8 (.D(data[7]), .CK(mem_22__7__N_174), .Q(\mem[22] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5067_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i2 (.D(data[1]), .CK(mem_21__7__N_171), .Q(\mem[21] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i3 (.D(data[2]), .CK(mem_21__7__N_171), .Q(\mem[21] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i4 (.D(data[3]), .CK(mem_21__7__N_171), .Q(\mem[21] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i5 (.D(data[4]), .CK(mem_21__7__N_171), .Q(\mem[21] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i6 (.D(data[5]), .CK(mem_21__7__N_171), .Q(\mem[21] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i7 (.D(data[6]), .CK(mem_21__7__N_171), .Q(\mem[21] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5064_i8 (.D(data[7]), .CK(mem_21__7__N_171), .Q(\mem[21] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5064_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5061_i2 (.D(data[1]), .CK(mem_20__7__N_168), .Q(\mem[20] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5061_i3 (.D(data[2]), .CK(mem_20__7__N_168), .Q(\mem[20] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5061_i4 (.D(data[3]), .CK(mem_20__7__N_168), .Q(\mem[20] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5061_i5 (.D(data[4]), .CK(mem_20__7__N_168), .Q(\mem[20] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5061_i6 (.D(data[5]), .CK(mem_20__7__N_168), .Q(\mem[20] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5061_i7 (.D(data[6]), .CK(mem_20__7__N_168), .Q(\mem[20] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5061_i8 (.D(data[7]), .CK(mem_20__7__N_168), .Q(\mem[20] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5061_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i2 (.D(data[1]), .CK(mem_19__7__N_165), .Q(\mem[19] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i3 (.D(data[2]), .CK(mem_19__7__N_165), .Q(\mem[19] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i4 (.D(data[3]), .CK(mem_19__7__N_165), .Q(\mem[19] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i5 (.D(data[4]), .CK(mem_19__7__N_165), .Q(\mem[19] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i6 (.D(data[5]), .CK(mem_19__7__N_165), .Q(\mem[19] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i7 (.D(data[6]), .CK(mem_19__7__N_165), .Q(\mem[19] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5058_i8 (.D(data[7]), .CK(mem_19__7__N_165), .Q(\mem[19] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5058_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5055_i2 (.D(data[1]), .CK(mem_18__7__N_162), .Q(\mem[18] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5055_i3 (.D(data[2]), .CK(mem_18__7__N_162), .Q(\mem[18] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5055_i4 (.D(data[3]), .CK(mem_18__7__N_162), .Q(\mem[18] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5055_i5 (.D(data[4]), .CK(mem_18__7__N_162), .Q(\mem[18] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5055_i6 (.D(data[5]), .CK(mem_18__7__N_162), .Q(\mem[18] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5055_i7 (.D(data[6]), .CK(mem_18__7__N_162), .Q(\mem[18] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5055_i8 (.D(data[7]), .CK(mem_18__7__N_162), .Q(\mem[18] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5055_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5052_i2 (.D(data[1]), .CK(mem_17__7__N_159), .Q(\mem[17] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5052_i3 (.D(data[2]), .CK(mem_17__7__N_159), .Q(\mem[17] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5052_i4 (.D(data[3]), .CK(mem_17__7__N_159), .Q(\mem[17] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5052_i5 (.D(data[4]), .CK(mem_17__7__N_159), .Q(\mem[17] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5052_i6 (.D(data[5]), .CK(mem_17__7__N_159), .Q(\mem[17] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5052_i7 (.D(data[6]), .CK(mem_17__7__N_159), .Q(\mem[17] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5052_i8 (.D(data[7]), .CK(mem_17__7__N_159), .Q(\mem[17] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5052_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i2 (.D(data[1]), .CK(mem_16__7__N_156), .Q(\mem[16] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i3 (.D(data[2]), .CK(mem_16__7__N_156), .Q(\mem[16] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i4 (.D(data[3]), .CK(mem_16__7__N_156), .Q(\mem[16] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i5 (.D(data[4]), .CK(mem_16__7__N_156), .Q(\mem[16] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i6 (.D(data[5]), .CK(mem_16__7__N_156), .Q(\mem[16] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i7 (.D(data[6]), .CK(mem_16__7__N_156), .Q(\mem[16] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5049_i8 (.D(data[7]), .CK(mem_16__7__N_156), .Q(\mem[16] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5049_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5046_i2 (.D(data[1]), .CK(mem_15__7__N_153), .Q(\mem[15] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5046_i3 (.D(data[2]), .CK(mem_15__7__N_153), .Q(\mem[15] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5046_i4 (.D(data[3]), .CK(mem_15__7__N_153), .Q(\mem[15] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5046_i5 (.D(data[4]), .CK(mem_15__7__N_153), .Q(\mem[15] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5046_i6 (.D(data[5]), .CK(mem_15__7__N_153), .Q(\mem[15] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5046_i7 (.D(data[6]), .CK(mem_15__7__N_153), .Q(\mem[15] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5046_i8 (.D(data[7]), .CK(mem_15__7__N_153), .Q(\mem[15] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5046_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5043_i2 (.D(data[1]), .CK(mem_14__7__N_150), .Q(\mem[14] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5043_i3 (.D(data[2]), .CK(mem_14__7__N_150), .Q(\mem[14] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5043_i4 (.D(data[3]), .CK(mem_14__7__N_150), .Q(\mem[14] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5043_i5 (.D(data[4]), .CK(mem_14__7__N_150), .Q(\mem[14] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5043_i6 (.D(data[5]), .CK(mem_14__7__N_150), .Q(\mem[14] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5043_i7 (.D(data[6]), .CK(mem_14__7__N_150), .Q(\mem[14] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5043_i8 (.D(data[7]), .CK(mem_14__7__N_150), .Q(\mem[14] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5043_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5040_i2 (.D(data[1]), .CK(mem_13__7__N_147), .Q(\mem[13] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5040_i3 (.D(data[2]), .CK(mem_13__7__N_147), .Q(\mem[13] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5040_i4 (.D(data[3]), .CK(mem_13__7__N_147), .Q(\mem[13] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5040_i5 (.D(data[4]), .CK(mem_13__7__N_147), .Q(\mem[13] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5040_i6 (.D(data[5]), .CK(mem_13__7__N_147), .Q(\mem[13] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5040_i7 (.D(data[6]), .CK(mem_13__7__N_147), .Q(\mem[13] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5040_i8 (.D(data[7]), .CK(mem_13__7__N_147), .Q(\mem[13] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5040_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5037_i2 (.D(data[1]), .CK(mem_12__7__N_144), .Q(\mem[12] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5037_i3 (.D(data[2]), .CK(mem_12__7__N_144), .Q(\mem[12] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5037_i4 (.D(data[3]), .CK(mem_12__7__N_144), .Q(\mem[12] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5037_i5 (.D(data[4]), .CK(mem_12__7__N_144), .Q(\mem[12] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5037_i6 (.D(data[5]), .CK(mem_12__7__N_144), .Q(\mem[12] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5037_i7 (.D(data[6]), .CK(mem_12__7__N_144), .Q(\mem[12] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5037_i8 (.D(data[7]), .CK(mem_12__7__N_144), .Q(\mem[12] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5037_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i2 (.D(data[1]), .CK(mem_11__7__N_141), .Q(\mem[11] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i3 (.D(data[2]), .CK(mem_11__7__N_141), .Q(\mem[11] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i4 (.D(data[3]), .CK(mem_11__7__N_141), .Q(\mem[11] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i5 (.D(data[4]), .CK(mem_11__7__N_141), .Q(\mem[11] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i6 (.D(data[5]), .CK(mem_11__7__N_141), .Q(\mem[11] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i7 (.D(data[6]), .CK(mem_11__7__N_141), .Q(\mem[11] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5034_i8 (.D(data[7]), .CK(mem_11__7__N_141), .Q(\mem[11] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5034_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5031_i2 (.D(data[1]), .CK(mem_10__7__N_138), .Q(\mem[10] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5031_i3 (.D(data[2]), .CK(mem_10__7__N_138), .Q(\mem[10] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5031_i4 (.D(data[3]), .CK(mem_10__7__N_138), .Q(\mem[10] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5031_i5 (.D(data[4]), .CK(mem_10__7__N_138), .Q(\mem[10] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5031_i6 (.D(data[5]), .CK(mem_10__7__N_138), .Q(\mem[10] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5031_i7 (.D(data[6]), .CK(mem_10__7__N_138), .Q(\mem[10] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5031_i8 (.D(data[7]), .CK(mem_10__7__N_138), .Q(\mem[10] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5031_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5028_i2 (.D(data[1]), .CK(mem_9__7__N_135), .Q(\mem[9] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5028_i3 (.D(data[2]), .CK(mem_9__7__N_135), .Q(\mem[9] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5028_i4 (.D(data[3]), .CK(mem_9__7__N_135), .Q(\mem[9] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5028_i5 (.D(data[4]), .CK(mem_9__7__N_135), .Q(\mem[9] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5028_i6 (.D(data[5]), .CK(mem_9__7__N_135), .Q(\mem[9] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5028_i7 (.D(data[6]), .CK(mem_9__7__N_135), .Q(\mem[9] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5028_i8 (.D(data[7]), .CK(mem_9__7__N_135), .Q(\mem[9] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5028_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5025_i2 (.D(data[1]), .CK(mem_8__7__N_132), .Q(\mem[8] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5025_i3 (.D(data[2]), .CK(mem_8__7__N_132), .Q(\mem[8] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5025_i4 (.D(data[3]), .CK(mem_8__7__N_132), .Q(\mem[8] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5025_i5 (.D(data[4]), .CK(mem_8__7__N_132), .Q(\mem[8] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5025_i6 (.D(data[5]), .CK(mem_8__7__N_132), .Q(\mem[8] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5025_i7 (.D(data[6]), .CK(mem_8__7__N_132), .Q(\mem[8] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5025_i8 (.D(data[7]), .CK(mem_8__7__N_132), .Q(\mem[8] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5025_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5022_i2 (.D(data[1]), .CK(mem_7__7__N_129), .Q(\mem[7] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5022_i3 (.D(data[2]), .CK(mem_7__7__N_129), .Q(\mem[7] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5022_i4 (.D(data[3]), .CK(mem_7__7__N_129), .Q(\mem[7] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5022_i5 (.D(data[4]), .CK(mem_7__7__N_129), .Q(\mem[7] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5022_i6 (.D(data[5]), .CK(mem_7__7__N_129), .Q(\mem[7] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5022_i7 (.D(data[6]), .CK(mem_7__7__N_129), .Q(\mem[7] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5022_i8 (.D(data[7]), .CK(mem_7__7__N_129), .Q(\mem[7] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5022_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5019_i2 (.D(data[1]), .CK(mem_6__7__N_126), .Q(\mem[6] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5019_i3 (.D(data[2]), .CK(mem_6__7__N_126), .Q(\mem[6] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5019_i4 (.D(data[3]), .CK(mem_6__7__N_126), .Q(\mem[6] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5019_i5 (.D(data[4]), .CK(mem_6__7__N_126), .Q(\mem[6] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5019_i6 (.D(data[5]), .CK(mem_6__7__N_126), .Q(\mem[6] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5019_i7 (.D(data[6]), .CK(mem_6__7__N_126), .Q(\mem[6] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5019_i8 (.D(data[7]), .CK(mem_6__7__N_126), .Q(\mem[6] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5019_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5016_i2 (.D(data[1]), .CK(mem_5__7__N_123), .Q(\mem[5] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5016_i3 (.D(data[2]), .CK(mem_5__7__N_123), .Q(\mem[5] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5016_i4 (.D(data[3]), .CK(mem_5__7__N_123), .Q(\mem[5] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5016_i5 (.D(data[4]), .CK(mem_5__7__N_123), .Q(\mem[5] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5016_i6 (.D(data[5]), .CK(mem_5__7__N_123), .Q(\mem[5] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5016_i7 (.D(data[6]), .CK(mem_5__7__N_123), .Q(\mem[5] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5016_i8 (.D(data[7]), .CK(mem_5__7__N_123), .Q(\mem[5] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5016_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5013_i2 (.D(data[1]), .CK(mem_4__7__N_120), .Q(\mem[4] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5013_i3 (.D(data[2]), .CK(mem_4__7__N_120), .Q(\mem[4] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5013_i4 (.D(data[3]), .CK(mem_4__7__N_120), .Q(\mem[4] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5013_i5 (.D(data[4]), .CK(mem_4__7__N_120), .Q(\mem[4] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5013_i6 (.D(data[5]), .CK(mem_4__7__N_120), .Q(\mem[4] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5013_i7 (.D(data[6]), .CK(mem_4__7__N_120), .Q(\mem[4] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5013_i8 (.D(data[7]), .CK(mem_4__7__N_120), .Q(\mem[4] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5013_i8.GSR = "DISABLED";
    FD1S1A data_7__I_0_5010_i2 (.D(data[1]), .CK(mem_3__7__N_117), .Q(\mem[3] [1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i2.GSR = "DISABLED";
    FD1S1A data_7__I_0_5010_i3 (.D(data[2]), .CK(mem_3__7__N_117), .Q(\mem[3] [2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i3.GSR = "DISABLED";
    FD1S1A data_7__I_0_5010_i4 (.D(data[3]), .CK(mem_3__7__N_117), .Q(\mem[3] [3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i4.GSR = "DISABLED";
    FD1S1A data_7__I_0_5010_i5 (.D(data[4]), .CK(mem_3__7__N_117), .Q(\mem[3] [4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i5.GSR = "DISABLED";
    FD1S1A data_7__I_0_5010_i6 (.D(data[5]), .CK(mem_3__7__N_117), .Q(\mem[3] [5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i6.GSR = "DISABLED";
    FD1S1A data_7__I_0_5010_i7 (.D(data[6]), .CK(mem_3__7__N_117), .Q(\mem[3] [6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i7.GSR = "DISABLED";
    FD1S1A data_7__I_0_5010_i8 (.D(data[7]), .CK(mem_3__7__N_117), .Q(\mem[3] [7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=20, LSE_LCOL=10, LSE_RCOL=19, LSE_LLINE=44, LSE_RLINE=44 */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(59[2] 83[14])
    defparam data_7__I_0_5010_i8.GSR = "DISABLED";
    PFUMX i2458032_i1 (.BLUT(n44436), .ALUT(n44467), .C0(address[5]), 
          .Z(data_7__N_89[5]));
    PFUMX i2457429_i1 (.BLUT(n44405), .ALUT(n44498), .C0(address[5]), 
          .Z(data_7__N_89[4]));
    PFUMX i2456826_i1 (.BLUT(n44374), .ALUT(n44529), .C0(address[5]), 
          .Z(data_7__N_89[3]));
    PFUMX i2456223_i1 (.BLUT(n44343), .ALUT(n44560), .C0(address[5]), 
          .Z(data_7__N_89[2]));
    PFUMX i2455620_i1 (.BLUT(n44312), .ALUT(n44591), .C0(address[5]), 
          .Z(data_7__N_89[1]));
    PFUMX i2455017_i1 (.BLUT(n44281), .ALUT(n44622), .C0(address[5]), 
          .Z(data_7__N_89[0]));
    PFUMX i2454414_i1 (.BLUT(n44250), .ALUT(n44653), .C0(address[5]), 
          .Z(data_7__N_89[7]));
    PFUMX i2453811_i1 (.BLUT(n44219), .ALUT(n44684), .C0(address[5]), 
          .Z(data_7__N_89[6]));
    L6MUX21 i37725 (.D0(n44616), .D1(n44617), .SD(address[3]), .Z(n44620));
    L6MUX21 i37726 (.D0(n44618), .D1(n44619), .SD(address[3]), .Z(n44621));
    L6MUX21 i37756 (.D0(n44647), .D1(n44648), .SD(address[3]), .Z(n44651));
    L6MUX21 i37757 (.D0(n44649), .D1(n44650), .SD(address[3]), .Z(n44652));
    L6MUX21 i37787 (.D0(n44678), .D1(n44679), .SD(address[3]), .Z(n44682));
    L6MUX21 i37788 (.D0(n44680), .D1(n44681), .SD(address[3]), .Z(n44683));
    L6MUX21 i37322 (.D0(n44213), .D1(n44214), .SD(address[3]), .Z(n44217));
    L6MUX21 i37323 (.D0(n44215), .D1(n44216), .SD(address[3]), .Z(n44218));
    L6MUX21 i37353 (.D0(n44244), .D1(n44245), .SD(address[3]), .Z(n44248));
    L6MUX21 i37354 (.D0(n44246), .D1(n44247), .SD(address[3]), .Z(n44249));
    L6MUX21 i37384 (.D0(n44275), .D1(n44276), .SD(address[3]), .Z(n44279));
    L6MUX21 i37385 (.D0(n44277), .D1(n44278), .SD(address[3]), .Z(n44280));
    L6MUX21 i37601 (.D0(n44492), .D1(n44493), .SD(address[3]), .Z(n44496));
    L6MUX21 i37602 (.D0(n44494), .D1(n44495), .SD(address[3]), .Z(n44497));
    L6MUX21 i37415 (.D0(n44306), .D1(n44307), .SD(address[3]), .Z(n44310));
    L6MUX21 i37416 (.D0(n44308), .D1(n44309), .SD(address[3]), .Z(n44311));
    L6MUX21 i37632 (.D0(n44523), .D1(n44524), .SD(address[3]), .Z(n44527));
    L6MUX21 i37633 (.D0(n44525), .D1(n44526), .SD(address[3]), .Z(n44528));
    L6MUX21 i37446 (.D0(n44337), .D1(n44338), .SD(address[3]), .Z(n44341));
    L6MUX21 i37447 (.D0(n44339), .D1(n44340), .SD(address[3]), .Z(n44342));
    L6MUX21 i37663 (.D0(n44554), .D1(n44555), .SD(address[3]), .Z(n44558));
    L6MUX21 i37664 (.D0(n44556), .D1(n44557), .SD(address[3]), .Z(n44559));
    L6MUX21 i37477 (.D0(n44368), .D1(n44369), .SD(address[3]), .Z(n44372));
    L6MUX21 i37478 (.D0(n44370), .D1(n44371), .SD(address[3]), .Z(n44373));
    L6MUX21 i37508 (.D0(n44399), .D1(n44400), .SD(address[3]), .Z(n44403));
    L6MUX21 i37509 (.D0(n44401), .D1(n44402), .SD(address[3]), .Z(n44404));
    L6MUX21 i37694 (.D0(n44585), .D1(n44586), .SD(address[3]), .Z(n44589));
    L6MUX21 i37695 (.D0(n44587), .D1(n44588), .SD(address[3]), .Z(n44590));
    L6MUX21 i37539 (.D0(n44430), .D1(n44431), .SD(address[3]), .Z(n44434));
    L6MUX21 i37540 (.D0(n44432), .D1(n44433), .SD(address[3]), .Z(n44435));
    L6MUX21 i37570 (.D0(n44461), .D1(n44462), .SD(address[3]), .Z(n44465));
    L6MUX21 i37571 (.D0(n44463), .D1(n44464), .SD(address[3]), .Z(n44466));
    L6MUX21 i37721 (.D0(n44608), .D1(n44609), .SD(address[2]), .Z(n44616));
    L6MUX21 i37722 (.D0(n44610), .D1(n44611), .SD(address[2]), .Z(n44617));
    L6MUX21 i37723 (.D0(n44612), .D1(n44613), .SD(address[2]), .Z(n44618));
    L6MUX21 i37724 (.D0(n44614), .D1(n44615), .SD(address[2]), .Z(n44619));
    PFUMX i37563 (.BLUT(n44447), .ALUT(n44448), .C0(address[1]), .Z(n44458));
    L6MUX21 i37318 (.D0(n44205), .D1(n44206), .SD(address[2]), .Z(n44213));
    L6MUX21 i37752 (.D0(n44639), .D1(n44640), .SD(address[2]), .Z(n44647));
    L6MUX21 i37319 (.D0(n44207), .D1(n44208), .SD(address[2]), .Z(n44214));
    L6MUX21 i37753 (.D0(n44641), .D1(n44642), .SD(address[2]), .Z(n44648));
    L6MUX21 i37754 (.D0(n44643), .D1(n44644), .SD(address[2]), .Z(n44649));
    L6MUX21 i37755 (.D0(n44645), .D1(n44646), .SD(address[2]), .Z(n44650));
    L6MUX21 i37320 (.D0(n44209), .D1(n44210), .SD(address[2]), .Z(n44215));
    L6MUX21 i37783 (.D0(n44670), .D1(n44671), .SD(address[2]), .Z(n44678));
    L6MUX21 i37784 (.D0(n44672), .D1(n44673), .SD(address[2]), .Z(n44679));
    L6MUX21 i37785 (.D0(n44674), .D1(n44675), .SD(address[2]), .Z(n44680));
    L6MUX21 i37786 (.D0(n44676), .D1(n44677), .SD(address[2]), .Z(n44681));
    L6MUX21 i37321 (.D0(n44211), .D1(n44212), .SD(address[2]), .Z(n44216));
    L6MUX21 i37349 (.D0(n44236), .D1(n44237), .SD(address[2]), .Z(n44244));
    L6MUX21 i37350 (.D0(n44238), .D1(n44239), .SD(address[2]), .Z(n44245));
    L6MUX21 i37351 (.D0(n44240), .D1(n44241), .SD(address[2]), .Z(n44246));
    L6MUX21 i37352 (.D0(n44242), .D1(n44243), .SD(address[2]), .Z(n44247));
    L6MUX21 i37597 (.D0(n44484), .D1(n44485), .SD(address[2]), .Z(n44492));
    L6MUX21 i37598 (.D0(n44486), .D1(n44487), .SD(address[2]), .Z(n44493));
    L6MUX21 i37380 (.D0(n44267), .D1(n44268), .SD(address[2]), .Z(n44275));
    L6MUX21 i37381 (.D0(n44269), .D1(n44270), .SD(address[2]), .Z(n44276));
    L6MUX21 i37382 (.D0(n44271), .D1(n44272), .SD(address[2]), .Z(n44277));
    L6MUX21 i37383 (.D0(n44273), .D1(n44274), .SD(address[2]), .Z(n44278));
    L6MUX21 i37599 (.D0(n44488), .D1(n44489), .SD(address[2]), .Z(n44494));
    L6MUX21 i37600 (.D0(n44490), .D1(n44491), .SD(address[2]), .Z(n44495));
    L6MUX21 i37411 (.D0(n44298), .D1(n44299), .SD(address[2]), .Z(n44306));
    L6MUX21 i37412 (.D0(n44300), .D1(n44301), .SD(address[2]), .Z(n44307));
    L6MUX21 i37413 (.D0(n44302), .D1(n44303), .SD(address[2]), .Z(n44308));
    L6MUX21 i37414 (.D0(n44304), .D1(n44305), .SD(address[2]), .Z(n44309));
    L6MUX21 i37628 (.D0(n44515), .D1(n44516), .SD(address[2]), .Z(n44523));
    L6MUX21 i37629 (.D0(n44517), .D1(n44518), .SD(address[2]), .Z(n44524));
    L6MUX21 i37630 (.D0(n44519), .D1(n44520), .SD(address[2]), .Z(n44525));
    L6MUX21 i37631 (.D0(n44521), .D1(n44522), .SD(address[2]), .Z(n44526));
    L6MUX21 i37442 (.D0(n44329), .D1(n44330), .SD(address[2]), .Z(n44337));
    L6MUX21 i37443 (.D0(n44331), .D1(n44332), .SD(address[2]), .Z(n44338));
    L6MUX21 i37444 (.D0(n44333), .D1(n44334), .SD(address[2]), .Z(n44339));
    L6MUX21 i37445 (.D0(n44335), .D1(n44336), .SD(address[2]), .Z(n44340));
    L6MUX21 i37659 (.D0(n44546), .D1(n44547), .SD(address[2]), .Z(n44554));
    L6MUX21 i37660 (.D0(n44548), .D1(n44549), .SD(address[2]), .Z(n44555));
    L6MUX21 i37661 (.D0(n44550), .D1(n44551), .SD(address[2]), .Z(n44556));
    L6MUX21 i37662 (.D0(n44552), .D1(n44553), .SD(address[2]), .Z(n44557));
    L6MUX21 i37473 (.D0(n44360), .D1(n44361), .SD(address[2]), .Z(n44368));
    L6MUX21 i37474 (.D0(n44362), .D1(n44363), .SD(address[2]), .Z(n44369));
    L6MUX21 i37475 (.D0(n44364), .D1(n44365), .SD(address[2]), .Z(n44370));
    L6MUX21 i37476 (.D0(n44366), .D1(n44367), .SD(address[2]), .Z(n44371));
    L6MUX21 i37504 (.D0(n44391), .D1(n44392), .SD(address[2]), .Z(n44399));
    L6MUX21 i37505 (.D0(n44393), .D1(n44394), .SD(address[2]), .Z(n44400));
    L6MUX21 i37506 (.D0(n44395), .D1(n44396), .SD(address[2]), .Z(n44401));
    L6MUX21 i37507 (.D0(n44397), .D1(n44398), .SD(address[2]), .Z(n44402));
    L6MUX21 i37690 (.D0(n44577), .D1(n44578), .SD(address[2]), .Z(n44585));
    L6MUX21 i37691 (.D0(n44579), .D1(n44580), .SD(address[2]), .Z(n44586));
    L6MUX21 i37692 (.D0(n44581), .D1(n44582), .SD(address[2]), .Z(n44587));
    L6MUX21 i37535 (.D0(n44422), .D1(n44423), .SD(address[2]), .Z(n44430));
    L6MUX21 i37693 (.D0(n44583), .D1(n44584), .SD(address[2]), .Z(n44588));
    L6MUX21 i37536 (.D0(n44424), .D1(n44425), .SD(address[2]), .Z(n44431));
    L6MUX21 i37537 (.D0(n44426), .D1(n44427), .SD(address[2]), .Z(n44432));
    L6MUX21 i37538 (.D0(n44428), .D1(n44429), .SD(address[2]), .Z(n44433));
    L6MUX21 i37566 (.D0(n44453), .D1(n44454), .SD(address[2]), .Z(n44461));
    L6MUX21 i37567 (.D0(n44455), .D1(n44456), .SD(address[2]), .Z(n44462));
    L6MUX21 i37568 (.D0(n44457), .D1(n44458), .SD(address[2]), .Z(n44463));
    L6MUX21 i37569 (.D0(n44459), .D1(n44460), .SD(address[2]), .Z(n44464));
    PFUMX i37310 (.BLUT(n44189), .ALUT(n44190), .C0(address[1]), .Z(n44205));
    LUT4 i1_2_lut_rep_1152 (.A(address[5]), .B(address[4]), .Z(n46273)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_rep_1152.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_1115_3_lut (.A(address[5]), .B(address[4]), .C(address[3]), 
         .Z(n46236)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_rep_1115_3_lut.init = 16'hfbfb;
    LUT4 i1_2_lut_rep_1117_3_lut (.A(address[5]), .B(address[4]), .C(address[3]), 
         .Z(n46238)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_rep_1117_3_lut.init = 16'hbfbf;
    PFUMX i37311 (.BLUT(n44191), .ALUT(n44192), .C0(address[1]), .Z(n44206));
    PFUMX i37564 (.BLUT(n44449), .ALUT(n44450), .C0(address[1]), .Z(n44459));
    PFUMX i37312 (.BLUT(n44193), .ALUT(n44194), .C0(address[1]), .Z(n44207));
    PFUMX i37313 (.BLUT(n44195), .ALUT(n44196), .C0(address[1]), .Z(n44208));
    PFUMX i37314 (.BLUT(n44197), .ALUT(n44198), .C0(address[1]), .Z(n44209));
    PFUMX i37315 (.BLUT(n44199), .ALUT(n44200), .C0(address[1]), .Z(n44210));
    PFUMX i37744 (.BLUT(n44623), .ALUT(n44624), .C0(address[1]), .Z(n44639));
    PFUMX i37316 (.BLUT(n44201), .ALUT(n44202), .C0(address[1]), .Z(n44211));
    PFUMX i37745 (.BLUT(n44625), .ALUT(n44626), .C0(address[1]), .Z(n44640));
    PFUMX i37317 (.BLUT(n44203), .ALUT(n44204), .C0(address[1]), .Z(n44212));
    PFUMX i37746 (.BLUT(n44627), .ALUT(n44628), .C0(address[1]), .Z(n44641));
    LUT4 i1_2_lut_rep_1153 (.A(address[4]), .B(address[3]), .Z(n46274)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_rep_1153.init = 16'heeee;
    PFUMX i37747 (.BLUT(n44629), .ALUT(n44630), .C0(address[1]), .Z(n44642));
    LUT4 i1_2_lut_rep_1111_3_lut (.A(address[4]), .B(address[3]), .C(address[5]), 
         .Z(n46232)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_rep_1111_3_lut.init = 16'hfefe;
    PFUMX i37748 (.BLUT(n44631), .ALUT(n44632), .C0(address[1]), .Z(n44643));
    PFUMX i37749 (.BLUT(n44633), .ALUT(n44634), .C0(address[1]), .Z(n44644));
    PFUMX i37750 (.BLUT(n44635), .ALUT(n44636), .C0(address[1]), .Z(n44645));
    PFUMX i37751 (.BLUT(n44637), .ALUT(n44638), .C0(address[1]), .Z(n44646));
    PFUMX i37775 (.BLUT(n44654), .ALUT(n44655), .C0(address[1]), .Z(n44670));
    PFUMX i37776 (.BLUT(n44656), .ALUT(n44657), .C0(address[1]), .Z(n44671));
    PFUMX i37777 (.BLUT(n44658), .ALUT(n44659), .C0(address[1]), .Z(n44672));
    PFUMX i37778 (.BLUT(n44660), .ALUT(n44661), .C0(address[1]), .Z(n44673));
    PFUMX i37779 (.BLUT(n44662), .ALUT(n44663), .C0(address[1]), .Z(n44674));
    PFUMX i37780 (.BLUT(n44664), .ALUT(n44665), .C0(address[1]), .Z(n44675));
    PFUMX i37781 (.BLUT(n44666), .ALUT(n44667), .C0(address[1]), .Z(n44676));
    PFUMX i37782 (.BLUT(n44668), .ALUT(n44669), .C0(address[1]), .Z(n44677));
    LUT4 i37712_3_lut (.A(\mem[62] [0]), .B(\mem[63] [0]), .C(address[0]), 
         .Z(n44607)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37712_3_lut.init = 16'hcaca;
    PFUMX i37341 (.BLUT(n44220), .ALUT(n44221), .C0(address[1]), .Z(n44236));
    PFUMX i37342 (.BLUT(n44222), .ALUT(n44223), .C0(address[1]), .Z(n44237));
    PFUMX i37343 (.BLUT(n44224), .ALUT(n44225), .C0(address[1]), .Z(n44238));
    PFUMX i37344 (.BLUT(n44226), .ALUT(n44227), .C0(address[1]), .Z(n44239));
    PFUMX i37345 (.BLUT(n44228), .ALUT(n44229), .C0(address[1]), .Z(n44240));
    PFUMX i37346 (.BLUT(n44230), .ALUT(n44231), .C0(address[1]), .Z(n44241));
    PFUMX i37347 (.BLUT(n44232), .ALUT(n44233), .C0(address[1]), .Z(n44242));
    PFUMX i37348 (.BLUT(n44234), .ALUT(n44235), .C0(address[1]), .Z(n44243));
    PFUMX i37589 (.BLUT(n44468), .ALUT(n44469), .C0(address[1]), .Z(n44484));
    LUT4 i37711_3_lut (.A(\mem[60] [0]), .B(\mem[61] [0]), .C(address[0]), 
         .Z(n44606)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37711_3_lut.init = 16'hcaca;
    PFUMX i37565 (.BLUT(n44451), .ALUT(n44452), .C0(address[1]), .Z(n44460));
    PFUMX i37590 (.BLUT(n44470), .ALUT(n44471), .C0(address[1]), .Z(n44485));
    PFUMX i37591 (.BLUT(n44472), .ALUT(n44473), .C0(address[1]), .Z(n44486));
    PFUMX i37592 (.BLUT(n44474), .ALUT(n44475), .C0(address[1]), .Z(n44487));
    LUT4 i37549_3_lut (.A(\mem[46] [5]), .B(\mem[47] [5]), .C(address[0]), 
         .Z(n44444)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37549_3_lut.init = 16'hcaca;
    LUT4 i37548_3_lut (.A(\mem[44] [5]), .B(\mem[45] [5]), .C(address[0]), 
         .Z(n44443)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37548_3_lut.init = 16'hcaca;
    LUT4 i37547_3_lut (.A(\mem[42] [5]), .B(\mem[43] [5]), .C(address[0]), 
         .Z(n44442)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37547_3_lut.init = 16'hcaca;
    LUT4 i37546_3_lut (.A(\mem[40] [5]), .B(\mem[41] [5]), .C(address[0]), 
         .Z(n44441)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37546_3_lut.init = 16'hcaca;
    LUT4 i37545_3_lut (.A(\mem[38] [5]), .B(\mem[39] [5]), .C(address[0]), 
         .Z(n44440)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37545_3_lut.init = 16'hcaca;
    LUT4 i37544_3_lut (.A(\mem[36] [5]), .B(\mem[37] [5]), .C(address[0]), 
         .Z(n44439)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37544_3_lut.init = 16'hcaca;
    PFUMX i37372 (.BLUT(n44251), .ALUT(n44252), .C0(address[1]), .Z(n44267));
    LUT4 i1_2_lut_rep_1118_3_lut (.A(address[4]), .B(address[3]), .C(address[5]), 
         .Z(n46239)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_rep_1118_3_lut.init = 16'hefef;
    LUT4 i37710_3_lut (.A(\mem[58] [0]), .B(\mem[59] [0]), .C(address[0]), 
         .Z(n44605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37710_3_lut.init = 16'hcaca;
    LUT4 i37709_3_lut (.A(\mem[56] [0]), .B(\mem[57] [0]), .C(address[0]), 
         .Z(n44604)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37709_3_lut.init = 16'hcaca;
    PFUMX i37373 (.BLUT(n44253), .ALUT(n44254), .C0(address[1]), .Z(n44268));
    LUT4 i37543_3_lut (.A(\mem[34] [5]), .B(\mem[35] [5]), .C(address[0]), 
         .Z(n44438)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37543_3_lut.init = 16'hcaca;
    LUT4 i37542_3_lut (.A(\mem[32] [5]), .B(\mem[33] [5]), .C(address[0]), 
         .Z(n44437)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37542_3_lut.init = 16'hcaca;
    LUT4 i37526_3_lut (.A(\mem[30] [5]), .B(\mem[31] [5]), .C(address[0]), 
         .Z(n44421)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37526_3_lut.init = 16'hcaca;
    LUT4 i37708_3_lut (.A(\mem[54] [0]), .B(\mem[55] [0]), .C(address[0]), 
         .Z(n44603)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37708_3_lut.init = 16'hcaca;
    LUT4 i37707_3_lut (.A(\mem[52] [0]), .B(\mem[53] [0]), .C(address[0]), 
         .Z(n44602)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37707_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_1154 (.A(address[4]), .B(address[3]), .Z(n46275)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_rep_1154.init = 16'hbbbb;
    PFUMX i37374 (.BLUT(n44255), .ALUT(n44256), .C0(address[1]), .Z(n44269));
    LUT4 i37525_3_lut (.A(\mem[28] [5]), .B(\mem[29] [5]), .C(address[0]), 
         .Z(n44420)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37525_3_lut.init = 16'hcaca;
    LUT4 i37524_3_lut (.A(\mem[26] [5]), .B(\mem[27] [5]), .C(address[0]), 
         .Z(n44419)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37524_3_lut.init = 16'hcaca;
    LUT4 i37523_3_lut (.A(\mem[24] [5]), .B(\mem[25] [5]), .C(address[0]), 
         .Z(n44418)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37523_3_lut.init = 16'hcaca;
    LUT4 i37522_3_lut (.A(\mem[22] [5]), .B(\mem[23] [5]), .C(address[0]), 
         .Z(n44417)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37522_3_lut.init = 16'hcaca;
    LUT4 i37521_3_lut (.A(\mem[20] [5]), .B(\mem[21] [5]), .C(address[0]), 
         .Z(n44416)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37521_3_lut.init = 16'hcaca;
    LUT4 i37520_3_lut (.A(\mem[18] [5]), .B(\mem[19] [5]), .C(address[0]), 
         .Z(n44415)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37520_3_lut.init = 16'hcaca;
    LUT4 i37519_3_lut (.A(\mem[16] [5]), .B(\mem[17] [5]), .C(address[0]), 
         .Z(n44414)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37519_3_lut.init = 16'hcaca;
    PFUMX i37593 (.BLUT(n44476), .ALUT(n44477), .C0(address[1]), .Z(n44488));
    LUT4 i37518_3_lut (.A(\mem[14] [5]), .B(\mem[15] [5]), .C(address[0]), 
         .Z(n44413)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37518_3_lut.init = 16'hcaca;
    LUT4 i37706_3_lut (.A(\mem[50] [0]), .B(\mem[51] [0]), .C(address[0]), 
         .Z(n44601)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37706_3_lut.init = 16'hcaca;
    LUT4 i37517_3_lut (.A(\mem[12] [5]), .B(\mem[13] [5]), .C(address[0]), 
         .Z(n44412)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37517_3_lut.init = 16'hcaca;
    LUT4 i37705_3_lut (.A(\mem[48] [0]), .B(\mem[49] [0]), .C(address[0]), 
         .Z(n44600)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37705_3_lut.init = 16'hcaca;
    LUT4 i37681_3_lut (.A(\mem[62] [1]), .B(\mem[63] [1]), .C(address[0]), 
         .Z(n44576)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37681_3_lut.init = 16'hcaca;
    LUT4 i37680_3_lut (.A(\mem[60] [1]), .B(\mem[61] [1]), .C(address[0]), 
         .Z(n44575)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37680_3_lut.init = 16'hcaca;
    LUT4 i37516_3_lut (.A(\mem[10] [5]), .B(\mem[11] [5]), .C(address[0]), 
         .Z(n44411)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37516_3_lut.init = 16'hcaca;
    LUT4 i37515_3_lut (.A(\mem[8] [5]), .B(\mem[9] [5]), .C(address[0]), 
         .Z(n44410)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37515_3_lut.init = 16'hcaca;
    LUT4 i37514_3_lut (.A(\mem[6] [5]), .B(\mem[7] [5]), .C(address[0]), 
         .Z(n44409)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37514_3_lut.init = 16'hcaca;
    LUT4 i37513_3_lut (.A(\mem[4] [5]), .B(\mem[5] [5]), .C(address[0]), 
         .Z(n44408)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37513_3_lut.init = 16'hcaca;
    PFUMX i37594 (.BLUT(n44478), .ALUT(n44479), .C0(address[1]), .Z(n44489));
    LUT4 i37512_3_lut (.A(\mem[2] [5]), .B(\mem[3] [5]), .C(address[0]), 
         .Z(n44407)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37512_3_lut.init = 16'hcaca;
    LUT4 i37511_3_lut (.A(\mem[0] [5]), .B(\mem[1] [5]), .C(address[0]), 
         .Z(n44406)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37511_3_lut.init = 16'hcaca;
    LUT4 i37679_3_lut (.A(\mem[58] [1]), .B(\mem[59] [1]), .C(address[0]), 
         .Z(n44574)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37679_3_lut.init = 16'hcaca;
    PFUMX i37595 (.BLUT(n44480), .ALUT(n44481), .C0(address[1]), .Z(n44490));
    LUT4 i37678_3_lut (.A(\mem[56] [1]), .B(\mem[57] [1]), .C(address[0]), 
         .Z(n44573)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37678_3_lut.init = 16'hcaca;
    LUT4 i37677_3_lut (.A(\mem[54] [1]), .B(\mem[55] [1]), .C(address[0]), 
         .Z(n44572)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37677_3_lut.init = 16'hcaca;
    PFUMX i37596 (.BLUT(n44482), .ALUT(n44483), .C0(address[1]), .Z(n44491));
    LUT4 i37676_3_lut (.A(\mem[52] [1]), .B(\mem[53] [1]), .C(address[0]), 
         .Z(n44571)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37676_3_lut.init = 16'hcaca;
    LUT4 i37675_3_lut (.A(\mem[50] [1]), .B(\mem[51] [1]), .C(address[0]), 
         .Z(n44570)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37675_3_lut.init = 16'hcaca;
    LUT4 i37674_3_lut (.A(\mem[48] [1]), .B(\mem[49] [1]), .C(address[0]), 
         .Z(n44569)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37674_3_lut.init = 16'hcaca;
    LUT4 i37673_3_lut (.A(\mem[46] [1]), .B(\mem[47] [1]), .C(address[0]), 
         .Z(n44568)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37673_3_lut.init = 16'hcaca;
    LUT4 i37672_3_lut (.A(\mem[44] [1]), .B(\mem[45] [1]), .C(address[0]), 
         .Z(n44567)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37672_3_lut.init = 16'hcaca;
    LUT4 i37671_3_lut (.A(\mem[42] [1]), .B(\mem[43] [1]), .C(address[0]), 
         .Z(n44566)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37671_3_lut.init = 16'hcaca;
    LUT4 i37670_3_lut (.A(\mem[40] [1]), .B(\mem[41] [1]), .C(address[0]), 
         .Z(n44565)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37670_3_lut.init = 16'hcaca;
    PFUMX i37375 (.BLUT(n44257), .ALUT(n44258), .C0(address[1]), .Z(n44270));
    LUT4 i37669_3_lut (.A(\mem[38] [1]), .B(\mem[39] [1]), .C(address[0]), 
         .Z(n44564)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37669_3_lut.init = 16'hcaca;
    LUT4 i37668_3_lut (.A(\mem[36] [1]), .B(\mem[37] [1]), .C(address[0]), 
         .Z(n44563)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37668_3_lut.init = 16'hcaca;
    LUT4 i37667_3_lut (.A(\mem[34] [1]), .B(\mem[35] [1]), .C(address[0]), 
         .Z(n44562)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37667_3_lut.init = 16'hcaca;
    LUT4 i37666_3_lut (.A(\mem[32] [1]), .B(\mem[33] [1]), .C(address[0]), 
         .Z(n44561)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37666_3_lut.init = 16'hcaca;
    LUT4 i37495_3_lut (.A(\mem[30] [4]), .B(\mem[31] [4]), .C(address[0]), 
         .Z(n44390)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37495_3_lut.init = 16'hcaca;
    LUT4 i37494_3_lut (.A(\mem[28] [4]), .B(\mem[29] [4]), .C(address[0]), 
         .Z(n44389)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37494_3_lut.init = 16'hcaca;
    LUT4 i37493_3_lut (.A(\mem[26] [4]), .B(\mem[27] [4]), .C(address[0]), 
         .Z(n44388)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37493_3_lut.init = 16'hcaca;
    LUT4 i37492_3_lut (.A(\mem[24] [4]), .B(\mem[25] [4]), .C(address[0]), 
         .Z(n44387)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37492_3_lut.init = 16'hcaca;
    LUT4 i37491_3_lut (.A(\mem[22] [4]), .B(\mem[23] [4]), .C(address[0]), 
         .Z(n44386)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37491_3_lut.init = 16'hcaca;
    LUT4 i37490_3_lut (.A(\mem[20] [4]), .B(\mem[21] [4]), .C(address[0]), 
         .Z(n44385)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37490_3_lut.init = 16'hcaca;
    LUT4 i37489_3_lut (.A(\mem[18] [4]), .B(\mem[19] [4]), .C(address[0]), 
         .Z(n44384)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37489_3_lut.init = 16'hcaca;
    LUT4 i37488_3_lut (.A(\mem[16] [4]), .B(\mem[17] [4]), .C(address[0]), 
         .Z(n44383)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37488_3_lut.init = 16'hcaca;
    PFUMX i37376 (.BLUT(n44259), .ALUT(n44260), .C0(address[1]), .Z(n44271));
    PFUMX i37377 (.BLUT(n44261), .ALUT(n44262), .C0(address[1]), .Z(n44272));
    LUT4 i37487_3_lut (.A(\mem[14] [4]), .B(\mem[15] [4]), .C(address[0]), 
         .Z(n44382)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37487_3_lut.init = 16'hcaca;
    PFUMX i37378 (.BLUT(n44263), .ALUT(n44264), .C0(address[1]), .Z(n44273));
    LUT4 i37486_3_lut (.A(\mem[12] [4]), .B(\mem[13] [4]), .C(address[0]), 
         .Z(n44381)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37486_3_lut.init = 16'hcaca;
    PFUMX i37713 (.BLUT(n44592), .ALUT(n44593), .C0(address[1]), .Z(n44608));
    LUT4 i37485_3_lut (.A(\mem[10] [4]), .B(\mem[11] [4]), .C(address[0]), 
         .Z(n44380)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37485_3_lut.init = 16'hcaca;
    LUT4 i37484_3_lut (.A(\mem[8] [4]), .B(\mem[9] [4]), .C(address[0]), 
         .Z(n44379)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37484_3_lut.init = 16'hcaca;
    LUT4 i37483_3_lut (.A(\mem[6] [4]), .B(\mem[7] [4]), .C(address[0]), 
         .Z(n44378)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37483_3_lut.init = 16'hcaca;
    PFUMX i37379 (.BLUT(n44265), .ALUT(n44266), .C0(address[1]), .Z(n44274));
    LUT4 i37482_3_lut (.A(\mem[4] [4]), .B(\mem[5] [4]), .C(address[0]), 
         .Z(n44377)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37482_3_lut.init = 16'hcaca;
    LUT4 i37481_3_lut (.A(\mem[2] [4]), .B(\mem[3] [4]), .C(address[0]), 
         .Z(n44376)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37481_3_lut.init = 16'hcaca;
    LUT4 i37480_3_lut (.A(\mem[0] [4]), .B(\mem[1] [4]), .C(address[0]), 
         .Z(n44375)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37480_3_lut.init = 16'hcaca;
    LUT4 i37464_3_lut (.A(\mem[30] [3]), .B(\mem[31] [3]), .C(address[0]), 
         .Z(n44359)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37464_3_lut.init = 16'hcaca;
    LUT4 i37463_3_lut (.A(\mem[28] [3]), .B(\mem[29] [3]), .C(address[0]), 
         .Z(n44358)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37463_3_lut.init = 16'hcaca;
    LUT4 i37462_3_lut (.A(\mem[26] [3]), .B(\mem[27] [3]), .C(address[0]), 
         .Z(n44357)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37462_3_lut.init = 16'hcaca;
    PFUMX i37620 (.BLUT(n44499), .ALUT(n44500), .C0(address[1]), .Z(n44515));
    LUT4 i37461_3_lut (.A(\mem[24] [3]), .B(\mem[25] [3]), .C(address[0]), 
         .Z(n44356)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37461_3_lut.init = 16'hcaca;
    LUT4 i37460_3_lut (.A(\mem[22] [3]), .B(\mem[23] [3]), .C(address[0]), 
         .Z(n44355)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37460_3_lut.init = 16'hcaca;
    LUT4 i37459_3_lut (.A(\mem[20] [3]), .B(\mem[21] [3]), .C(address[0]), 
         .Z(n44354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37459_3_lut.init = 16'hcaca;
    LUT4 i37458_3_lut (.A(\mem[18] [3]), .B(\mem[19] [3]), .C(address[0]), 
         .Z(n44353)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37458_3_lut.init = 16'hcaca;
    LUT4 i37457_3_lut (.A(\mem[16] [3]), .B(\mem[17] [3]), .C(address[0]), 
         .Z(n44352)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37457_3_lut.init = 16'hcaca;
    LUT4 i37456_3_lut (.A(\mem[14] [3]), .B(\mem[15] [3]), .C(address[0]), 
         .Z(n44351)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37456_3_lut.init = 16'hcaca;
    LUT4 i37455_3_lut (.A(\mem[12] [3]), .B(\mem[13] [3]), .C(address[0]), 
         .Z(n44350)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37455_3_lut.init = 16'hcaca;
    LUT4 i37454_3_lut (.A(\mem[10] [3]), .B(\mem[11] [3]), .C(address[0]), 
         .Z(n44349)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37454_3_lut.init = 16'hcaca;
    LUT4 i37453_3_lut (.A(\mem[8] [3]), .B(\mem[9] [3]), .C(address[0]), 
         .Z(n44348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37453_3_lut.init = 16'hcaca;
    LUT4 i37452_3_lut (.A(\mem[6] [3]), .B(\mem[7] [3]), .C(address[0]), 
         .Z(n44347)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37452_3_lut.init = 16'hcaca;
    LUT4 i37451_3_lut (.A(\mem[4] [3]), .B(\mem[5] [3]), .C(address[0]), 
         .Z(n44346)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37451_3_lut.init = 16'hcaca;
    PFUMX i37403 (.BLUT(n44282), .ALUT(n44283), .C0(address[1]), .Z(n44298));
    LUT4 i37450_3_lut (.A(\mem[2] [3]), .B(\mem[3] [3]), .C(address[0]), 
         .Z(n44345)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37450_3_lut.init = 16'hcaca;
    LUT4 i37449_3_lut (.A(\mem[0] [3]), .B(\mem[1] [3]), .C(address[0]), 
         .Z(n44344)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37449_3_lut.init = 16'hcaca;
    LUT4 i37650_3_lut (.A(\mem[62] [2]), .B(\mem[63] [2]), .C(address[0]), 
         .Z(n44545)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37650_3_lut.init = 16'hcaca;
    LUT4 i37649_3_lut (.A(\mem[60] [2]), .B(\mem[61] [2]), .C(address[0]), 
         .Z(n44544)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37649_3_lut.init = 16'hcaca;
    PFUMX i37404 (.BLUT(n44284), .ALUT(n44285), .C0(address[1]), .Z(n44299));
    PFUMX i37621 (.BLUT(n44501), .ALUT(n44502), .C0(address[1]), .Z(n44516));
    LUT4 i37648_3_lut (.A(\mem[58] [2]), .B(\mem[59] [2]), .C(address[0]), 
         .Z(n44543)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37648_3_lut.init = 16'hcaca;
    LUT4 i37647_3_lut (.A(\mem[56] [2]), .B(\mem[57] [2]), .C(address[0]), 
         .Z(n44542)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37647_3_lut.init = 16'hcaca;
    LUT4 i37646_3_lut (.A(\mem[54] [2]), .B(\mem[55] [2]), .C(address[0]), 
         .Z(n44541)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37646_3_lut.init = 16'hcaca;
    PFUMX i37405 (.BLUT(n44286), .ALUT(n44287), .C0(address[1]), .Z(n44300));
    LUT4 i37704_3_lut (.A(\mem[46] [0]), .B(\mem[47] [0]), .C(address[0]), 
         .Z(n44599)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37704_3_lut.init = 16'hcaca;
    LUT4 i37645_3_lut (.A(\mem[52] [2]), .B(\mem[53] [2]), .C(address[0]), 
         .Z(n44540)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37645_3_lut.init = 16'hcaca;
    LUT4 i37644_3_lut (.A(\mem[50] [2]), .B(\mem[51] [2]), .C(address[0]), 
         .Z(n44539)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37644_3_lut.init = 16'hcaca;
    LUT4 i37643_3_lut (.A(\mem[48] [2]), .B(\mem[49] [2]), .C(address[0]), 
         .Z(n44538)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37643_3_lut.init = 16'hcaca;
    LUT4 i37642_3_lut (.A(\mem[46] [2]), .B(\mem[47] [2]), .C(address[0]), 
         .Z(n44537)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37642_3_lut.init = 16'hcaca;
    LUT4 i37641_3_lut (.A(\mem[44] [2]), .B(\mem[45] [2]), .C(address[0]), 
         .Z(n44536)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37641_3_lut.init = 16'hcaca;
    LUT4 i37703_3_lut (.A(\mem[44] [0]), .B(\mem[45] [0]), .C(address[0]), 
         .Z(n44598)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37703_3_lut.init = 16'hcaca;
    LUT4 i37640_3_lut (.A(\mem[42] [2]), .B(\mem[43] [2]), .C(address[0]), 
         .Z(n44535)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37640_3_lut.init = 16'hcaca;
    LUT4 i37639_3_lut (.A(\mem[40] [2]), .B(\mem[41] [2]), .C(address[0]), 
         .Z(n44534)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37639_3_lut.init = 16'hcaca;
    LUT4 i37638_3_lut (.A(\mem[38] [2]), .B(\mem[39] [2]), .C(address[0]), 
         .Z(n44533)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37638_3_lut.init = 16'hcaca;
    LUT4 i37637_3_lut (.A(\mem[36] [2]), .B(\mem[37] [2]), .C(address[0]), 
         .Z(n44532)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37637_3_lut.init = 16'hcaca;
    LUT4 i37636_3_lut (.A(\mem[34] [2]), .B(\mem[35] [2]), .C(address[0]), 
         .Z(n44531)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37636_3_lut.init = 16'hcaca;
    LUT4 i37635_3_lut (.A(\mem[32] [2]), .B(\mem[33] [2]), .C(address[0]), 
         .Z(n44530)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37635_3_lut.init = 16'hcaca;
    LUT4 i37433_3_lut (.A(\mem[30] [2]), .B(\mem[31] [2]), .C(address[0]), 
         .Z(n44328)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37433_3_lut.init = 16'hcaca;
    LUT4 i37432_3_lut (.A(\mem[28] [2]), .B(\mem[29] [2]), .C(address[0]), 
         .Z(n44327)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37432_3_lut.init = 16'hcaca;
    LUT4 i37431_3_lut (.A(\mem[26] [2]), .B(\mem[27] [2]), .C(address[0]), 
         .Z(n44326)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37431_3_lut.init = 16'hcaca;
    LUT4 i37430_3_lut (.A(\mem[24] [2]), .B(\mem[25] [2]), .C(address[0]), 
         .Z(n44325)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37430_3_lut.init = 16'hcaca;
    PFUMX i37406 (.BLUT(n44288), .ALUT(n44289), .C0(address[1]), .Z(n44301));
    LUT4 i37429_3_lut (.A(\mem[22] [2]), .B(\mem[23] [2]), .C(address[0]), 
         .Z(n44324)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37429_3_lut.init = 16'hcaca;
    LUT4 i37428_3_lut (.A(\mem[20] [2]), .B(\mem[21] [2]), .C(address[0]), 
         .Z(n44323)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37428_3_lut.init = 16'hcaca;
    PFUMX i37407 (.BLUT(n44290), .ALUT(n44291), .C0(address[1]), .Z(n44302));
    LUT4 i37427_3_lut (.A(\mem[18] [2]), .B(\mem[19] [2]), .C(address[0]), 
         .Z(n44322)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37427_3_lut.init = 16'hcaca;
    LUT4 i37426_3_lut (.A(\mem[16] [2]), .B(\mem[17] [2]), .C(address[0]), 
         .Z(n44321)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37426_3_lut.init = 16'hcaca;
    LUT4 i37425_3_lut (.A(\mem[14] [2]), .B(\mem[15] [2]), .C(address[0]), 
         .Z(n44320)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37425_3_lut.init = 16'hcaca;
    LUT4 i37702_3_lut (.A(\mem[42] [0]), .B(\mem[43] [0]), .C(address[0]), 
         .Z(n44597)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37702_3_lut.init = 16'hcaca;
    LUT4 i37424_3_lut (.A(\mem[12] [2]), .B(\mem[13] [2]), .C(address[0]), 
         .Z(n44319)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37424_3_lut.init = 16'hcaca;
    PFUMX i37408 (.BLUT(n44292), .ALUT(n44293), .C0(address[1]), .Z(n44303));
    PFUMX i37714 (.BLUT(n44594), .ALUT(n44595), .C0(address[1]), .Z(n44609));
    PFUMX i37409 (.BLUT(n44294), .ALUT(n44295), .C0(address[1]), .Z(n44304));
    LUT4 i37423_3_lut (.A(\mem[10] [2]), .B(\mem[11] [2]), .C(address[0]), 
         .Z(n44318)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37423_3_lut.init = 16'hcaca;
    LUT4 i37422_3_lut (.A(\mem[8] [2]), .B(\mem[9] [2]), .C(address[0]), 
         .Z(n44317)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37422_3_lut.init = 16'hcaca;
    PFUMX i37410 (.BLUT(n44296), .ALUT(n44297), .C0(address[1]), .Z(n44305));
    PFUMX i37622 (.BLUT(n44503), .ALUT(n44504), .C0(address[1]), .Z(n44517));
    LUT4 i1_2_lut_rep_1113_3_lut (.A(address[4]), .B(address[3]), .C(address[5]), 
         .Z(n46234)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_rep_1113_3_lut.init = 16'hfbfb;
    LUT4 i37421_3_lut (.A(\mem[6] [2]), .B(\mem[7] [2]), .C(address[0]), 
         .Z(n44316)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37421_3_lut.init = 16'hcaca;
    LUT4 i37420_3_lut (.A(\mem[4] [2]), .B(\mem[5] [2]), .C(address[0]), 
         .Z(n44315)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37420_3_lut.init = 16'hcaca;
    LUT4 i37701_3_lut (.A(\mem[40] [0]), .B(\mem[41] [0]), .C(address[0]), 
         .Z(n44596)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37701_3_lut.init = 16'hcaca;
    LUT4 i37419_3_lut (.A(\mem[2] [2]), .B(\mem[3] [2]), .C(address[0]), 
         .Z(n44314)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37419_3_lut.init = 16'hcaca;
    PFUMX i37623 (.BLUT(n44505), .ALUT(n44506), .C0(address[1]), .Z(n44518));
    LUT4 i37418_3_lut (.A(\mem[0] [2]), .B(\mem[1] [2]), .C(address[0]), 
         .Z(n44313)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37418_3_lut.init = 16'hcaca;
    LUT4 i37619_3_lut (.A(\mem[62] [3]), .B(\mem[63] [3]), .C(address[0]), 
         .Z(n44514)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37619_3_lut.init = 16'hcaca;
    LUT4 i37618_3_lut (.A(\mem[60] [3]), .B(\mem[61] [3]), .C(address[0]), 
         .Z(n44513)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37618_3_lut.init = 16'hcaca;
    LUT4 i37617_3_lut (.A(\mem[58] [3]), .B(\mem[59] [3]), .C(address[0]), 
         .Z(n44512)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37617_3_lut.init = 16'hcaca;
    LUT4 i37616_3_lut (.A(\mem[56] [3]), .B(\mem[57] [3]), .C(address[0]), 
         .Z(n44511)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37616_3_lut.init = 16'hcaca;
    PFUMX i37624 (.BLUT(n44507), .ALUT(n44508), .C0(address[1]), .Z(n44519));
    LUT4 i37615_3_lut (.A(\mem[54] [3]), .B(\mem[55] [3]), .C(address[0]), 
         .Z(n44510)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37615_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_1120_3_lut (.A(address[4]), .B(address[3]), .C(address[5]), 
         .Z(n46241)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_rep_1120_3_lut.init = 16'hbfbf;
    PFUMX i37715 (.BLUT(n44596), .ALUT(n44597), .C0(address[1]), .Z(n44610));
    LUT4 i37614_3_lut (.A(\mem[52] [3]), .B(\mem[53] [3]), .C(address[0]), 
         .Z(n44509)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37614_3_lut.init = 16'hcaca;
    PFUMX i37625 (.BLUT(n44509), .ALUT(n44510), .C0(address[1]), .Z(n44520));
    LUT4 i37613_3_lut (.A(\mem[50] [3]), .B(\mem[51] [3]), .C(address[0]), 
         .Z(n44508)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37613_3_lut.init = 16'hcaca;
    PFUMX i37626 (.BLUT(n44511), .ALUT(n44512), .C0(address[1]), .Z(n44521));
    LUT4 i37612_3_lut (.A(\mem[48] [3]), .B(\mem[49] [3]), .C(address[0]), 
         .Z(n44507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37612_3_lut.init = 16'hcaca;
    LUT4 i37700_3_lut (.A(\mem[38] [0]), .B(\mem[39] [0]), .C(address[0]), 
         .Z(n44595)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37700_3_lut.init = 16'hcaca;
    LUT4 i37699_3_lut (.A(\mem[36] [0]), .B(\mem[37] [0]), .C(address[0]), 
         .Z(n44594)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37699_3_lut.init = 16'hcaca;
    LUT4 i37611_3_lut (.A(\mem[46] [3]), .B(\mem[47] [3]), .C(address[0]), 
         .Z(n44506)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37611_3_lut.init = 16'hcaca;
    LUT4 i37610_3_lut (.A(\mem[44] [3]), .B(\mem[45] [3]), .C(address[0]), 
         .Z(n44505)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37610_3_lut.init = 16'hcaca;
    LUT4 i37609_3_lut (.A(\mem[42] [3]), .B(\mem[43] [3]), .C(address[0]), 
         .Z(n44504)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37609_3_lut.init = 16'hcaca;
    LUT4 i37608_3_lut (.A(\mem[40] [3]), .B(\mem[41] [3]), .C(address[0]), 
         .Z(n44503)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37608_3_lut.init = 16'hcaca;
    PFUMX i37627 (.BLUT(n44513), .ALUT(n44514), .C0(address[1]), .Z(n44522));
    LUT4 i37402_3_lut (.A(\mem[30] [1]), .B(\mem[31] [1]), .C(address[0]), 
         .Z(n44297)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37402_3_lut.init = 16'hcaca;
    LUT4 i37401_3_lut (.A(\mem[28] [1]), .B(\mem[29] [1]), .C(address[0]), 
         .Z(n44296)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37401_3_lut.init = 16'hcaca;
    LUT4 i37400_3_lut (.A(\mem[26] [1]), .B(\mem[27] [1]), .C(address[0]), 
         .Z(n44295)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37400_3_lut.init = 16'hcaca;
    LUT4 i37399_3_lut (.A(\mem[24] [1]), .B(\mem[25] [1]), .C(address[0]), 
         .Z(n44294)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37399_3_lut.init = 16'hcaca;
    LUT4 i37398_3_lut (.A(\mem[22] [1]), .B(\mem[23] [1]), .C(address[0]), 
         .Z(n44293)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37398_3_lut.init = 16'hcaca;
    LUT4 i37397_3_lut (.A(\mem[20] [1]), .B(\mem[21] [1]), .C(address[0]), 
         .Z(n44292)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37397_3_lut.init = 16'hcaca;
    LUT4 i37396_3_lut (.A(\mem[18] [1]), .B(\mem[19] [1]), .C(address[0]), 
         .Z(n44291)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37396_3_lut.init = 16'hcaca;
    LUT4 i37395_3_lut (.A(\mem[16] [1]), .B(\mem[17] [1]), .C(address[0]), 
         .Z(n44290)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37395_3_lut.init = 16'hcaca;
    LUT4 i37394_3_lut (.A(\mem[14] [1]), .B(\mem[15] [1]), .C(address[0]), 
         .Z(n44289)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37394_3_lut.init = 16'hcaca;
    PFUMX i37434 (.BLUT(n44313), .ALUT(n44314), .C0(address[1]), .Z(n44329));
    LUT4 i37393_3_lut (.A(\mem[12] [1]), .B(\mem[13] [1]), .C(address[0]), 
         .Z(n44288)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37393_3_lut.init = 16'hcaca;
    PFUMX i37562 (.BLUT(n44445), .ALUT(n44446), .C0(address[1]), .Z(n44457));
    PFUMX i37435 (.BLUT(n44315), .ALUT(n44316), .C0(address[1]), .Z(n44330));
    LUT4 i37392_3_lut (.A(\mem[10] [1]), .B(\mem[11] [1]), .C(address[0]), 
         .Z(n44287)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37392_3_lut.init = 16'hcaca;
    LUT4 i37391_3_lut (.A(\mem[8] [1]), .B(\mem[9] [1]), .C(address[0]), 
         .Z(n44286)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37391_3_lut.init = 16'hcaca;
    LUT4 i37607_3_lut (.A(\mem[38] [3]), .B(\mem[39] [3]), .C(address[0]), 
         .Z(n44502)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37607_3_lut.init = 16'hcaca;
    LUT4 i37606_3_lut (.A(\mem[36] [3]), .B(\mem[37] [3]), .C(address[0]), 
         .Z(n44501)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37606_3_lut.init = 16'hcaca;
    LUT4 i37698_3_lut (.A(\mem[34] [0]), .B(\mem[35] [0]), .C(address[0]), 
         .Z(n44593)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37698_3_lut.init = 16'hcaca;
    LUT4 i37390_3_lut (.A(\mem[6] [1]), .B(\mem[7] [1]), .C(address[0]), 
         .Z(n44285)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37390_3_lut.init = 16'hcaca;
    LUT4 i37389_3_lut (.A(\mem[4] [1]), .B(\mem[5] [1]), .C(address[0]), 
         .Z(n44284)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37389_3_lut.init = 16'hcaca;
    PFUMX i37436 (.BLUT(n44317), .ALUT(n44318), .C0(address[1]), .Z(n44331));
    LUT4 i37388_3_lut (.A(\mem[2] [1]), .B(\mem[3] [1]), .C(address[0]), 
         .Z(n44283)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37388_3_lut.init = 16'hcaca;
    LUT4 i37387_3_lut (.A(\mem[0] [1]), .B(\mem[1] [1]), .C(address[0]), 
         .Z(n44282)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37387_3_lut.init = 16'hcaca;
    LUT4 i37605_3_lut (.A(\mem[34] [3]), .B(\mem[35] [3]), .C(address[0]), 
         .Z(n44500)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37605_3_lut.init = 16'hcaca;
    LUT4 i37604_3_lut (.A(\mem[32] [3]), .B(\mem[33] [3]), .C(address[0]), 
         .Z(n44499)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37604_3_lut.init = 16'hcaca;
    LUT4 i37697_3_lut (.A(\mem[32] [0]), .B(\mem[33] [0]), .C(address[0]), 
         .Z(n44592)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37697_3_lut.init = 16'hcaca;
    LUT4 i37371_3_lut (.A(\mem[30] [0]), .B(\mem[31] [0]), .C(address[0]), 
         .Z(n44266)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37371_3_lut.init = 16'hcaca;
    LUT4 i37370_3_lut (.A(\mem[28] [0]), .B(\mem[29] [0]), .C(address[0]), 
         .Z(n44265)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37370_3_lut.init = 16'hcaca;
    LUT4 i37369_3_lut (.A(\mem[26] [0]), .B(\mem[27] [0]), .C(address[0]), 
         .Z(n44264)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37369_3_lut.init = 16'hcaca;
    LUT4 i37368_3_lut (.A(\mem[24] [0]), .B(\mem[25] [0]), .C(address[0]), 
         .Z(n44263)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37368_3_lut.init = 16'hcaca;
    LUT4 i37367_3_lut (.A(\mem[22] [0]), .B(\mem[23] [0]), .C(address[0]), 
         .Z(n44262)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37367_3_lut.init = 16'hcaca;
    LUT4 i37366_3_lut (.A(\mem[20] [0]), .B(\mem[21] [0]), .C(address[0]), 
         .Z(n44261)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37366_3_lut.init = 16'hcaca;
    LUT4 i37365_3_lut (.A(\mem[18] [0]), .B(\mem[19] [0]), .C(address[0]), 
         .Z(n44260)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37365_3_lut.init = 16'hcaca;
    LUT4 i37364_3_lut (.A(\mem[16] [0]), .B(\mem[17] [0]), .C(address[0]), 
         .Z(n44259)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37364_3_lut.init = 16'hcaca;
    LUT4 i37363_3_lut (.A(\mem[14] [0]), .B(\mem[15] [0]), .C(address[0]), 
         .Z(n44258)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37363_3_lut.init = 16'hcaca;
    LUT4 i37557_3_lut (.A(\mem[62] [5]), .B(\mem[63] [5]), .C(address[0]), 
         .Z(n44452)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37557_3_lut.init = 16'hcaca;
    PFUMX i37437 (.BLUT(n44319), .ALUT(n44320), .C0(address[1]), .Z(n44332));
    LUT4 i37362_3_lut (.A(\mem[12] [0]), .B(\mem[13] [0]), .C(address[0]), 
         .Z(n44257)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37362_3_lut.init = 16'hcaca;
    LUT4 i37588_3_lut (.A(\mem[62] [4]), .B(\mem[63] [4]), .C(address[0]), 
         .Z(n44483)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37588_3_lut.init = 16'hcaca;
    LUT4 i37587_3_lut (.A(\mem[60] [4]), .B(\mem[61] [4]), .C(address[0]), 
         .Z(n44482)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37587_3_lut.init = 16'hcaca;
    LUT4 i37586_3_lut (.A(\mem[58] [4]), .B(\mem[59] [4]), .C(address[0]), 
         .Z(n44481)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37586_3_lut.init = 16'hcaca;
    LUT4 i37585_3_lut (.A(\mem[56] [4]), .B(\mem[57] [4]), .C(address[0]), 
         .Z(n44480)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37585_3_lut.init = 16'hcaca;
    LUT4 i37584_3_lut (.A(\mem[54] [4]), .B(\mem[55] [4]), .C(address[0]), 
         .Z(n44479)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37584_3_lut.init = 16'hcaca;
    LUT4 i37583_3_lut (.A(\mem[52] [4]), .B(\mem[53] [4]), .C(address[0]), 
         .Z(n44478)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37583_3_lut.init = 16'hcaca;
    LUT4 i37582_3_lut (.A(\mem[50] [4]), .B(\mem[51] [4]), .C(address[0]), 
         .Z(n44477)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37582_3_lut.init = 16'hcaca;
    PFUMX i37438 (.BLUT(n44321), .ALUT(n44322), .C0(address[1]), .Z(n44333));
    LUT4 i37581_3_lut (.A(\mem[48] [4]), .B(\mem[49] [4]), .C(address[0]), 
         .Z(n44476)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37581_3_lut.init = 16'hcaca;
    PFUMX i37439 (.BLUT(n44323), .ALUT(n44324), .C0(address[1]), .Z(n44334));
    LUT4 i37361_3_lut (.A(\mem[10] [0]), .B(\mem[11] [0]), .C(address[0]), 
         .Z(n44256)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37361_3_lut.init = 16'hcaca;
    PFUMX i37440 (.BLUT(n44325), .ALUT(n44326), .C0(address[1]), .Z(n44335));
    LUT4 i37360_3_lut (.A(\mem[8] [0]), .B(\mem[9] [0]), .C(address[0]), 
         .Z(n44255)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37360_3_lut.init = 16'hcaca;
    PFUMX i37441 (.BLUT(n44327), .ALUT(n44328), .C0(address[1]), .Z(n44336));
    LUT4 i37359_3_lut (.A(\mem[6] [0]), .B(\mem[7] [0]), .C(address[0]), 
         .Z(n44254)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37359_3_lut.init = 16'hcaca;
    LUT4 i37358_3_lut (.A(\mem[4] [0]), .B(\mem[5] [0]), .C(address[0]), 
         .Z(n44253)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37358_3_lut.init = 16'hcaca;
    PFUMX i37651 (.BLUT(n44530), .ALUT(n44531), .C0(address[1]), .Z(n44546));
    LUT4 i37357_3_lut (.A(\mem[2] [0]), .B(\mem[3] [0]), .C(address[0]), 
         .Z(n44252)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37357_3_lut.init = 16'hcaca;
    PFUMX i37652 (.BLUT(n44532), .ALUT(n44533), .C0(address[1]), .Z(n44547));
    LUT4 i37356_3_lut (.A(\mem[0] [0]), .B(\mem[1] [0]), .C(address[0]), 
         .Z(n44251)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37356_3_lut.init = 16'hcaca;
    LUT4 i37580_3_lut (.A(\mem[46] [4]), .B(\mem[47] [4]), .C(address[0]), 
         .Z(n44475)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37580_3_lut.init = 16'hcaca;
    LUT4 i37579_3_lut (.A(\mem[44] [4]), .B(\mem[45] [4]), .C(address[0]), 
         .Z(n44474)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37579_3_lut.init = 16'hcaca;
    PFUMX i37653 (.BLUT(n44534), .ALUT(n44535), .C0(address[1]), .Z(n44548));
    LUT4 i37578_3_lut (.A(\mem[42] [4]), .B(\mem[43] [4]), .C(address[0]), 
         .Z(n44473)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37578_3_lut.init = 16'hcaca;
    LUT4 i37577_3_lut (.A(\mem[40] [4]), .B(\mem[41] [4]), .C(address[0]), 
         .Z(n44472)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37577_3_lut.init = 16'hcaca;
    LUT4 i37576_3_lut (.A(\mem[38] [4]), .B(\mem[39] [4]), .C(address[0]), 
         .Z(n44471)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37576_3_lut.init = 16'hcaca;
    LUT4 i37575_3_lut (.A(\mem[36] [4]), .B(\mem[37] [4]), .C(address[0]), 
         .Z(n44470)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37575_3_lut.init = 16'hcaca;
    LUT4 i37556_3_lut (.A(\mem[60] [5]), .B(\mem[61] [5]), .C(address[0]), 
         .Z(n44451)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37556_3_lut.init = 16'hcaca;
    PFUMX i37716 (.BLUT(n44598), .ALUT(n44599), .C0(address[1]), .Z(n44611));
    PFUMX i37654 (.BLUT(n44536), .ALUT(n44537), .C0(address[1]), .Z(n44549));
    PFUMX i37655 (.BLUT(n44538), .ALUT(n44539), .C0(address[1]), .Z(n44550));
    LUT4 i37574_3_lut (.A(\mem[34] [4]), .B(\mem[35] [4]), .C(address[0]), 
         .Z(n44469)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37574_3_lut.init = 16'hcaca;
    PFUMX i37656 (.BLUT(n44540), .ALUT(n44541), .C0(address[1]), .Z(n44551));
    LUT4 i37573_3_lut (.A(\mem[32] [4]), .B(\mem[33] [4]), .C(address[0]), 
         .Z(n44468)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37573_3_lut.init = 16'hcaca;
    LUT4 i37340_3_lut (.A(\mem[30] [7]), .B(\mem[31] [7]), .C(address[0]), 
         .Z(n44235)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37340_3_lut.init = 16'hcaca;
    LUT4 i37339_3_lut (.A(\mem[28] [7]), .B(\mem[29] [7]), .C(address[0]), 
         .Z(n44234)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37339_3_lut.init = 16'hcaca;
    LUT4 i37338_3_lut (.A(\mem[26] [7]), .B(\mem[27] [7]), .C(address[0]), 
         .Z(n44233)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37338_3_lut.init = 16'hcaca;
    LUT4 i37337_3_lut (.A(\mem[24] [7]), .B(\mem[25] [7]), .C(address[0]), 
         .Z(n44232)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37337_3_lut.init = 16'hcaca;
    LUT4 i37336_3_lut (.A(\mem[22] [7]), .B(\mem[23] [7]), .C(address[0]), 
         .Z(n44231)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37336_3_lut.init = 16'hcaca;
    LUT4 i37335_3_lut (.A(\mem[20] [7]), .B(\mem[21] [7]), .C(address[0]), 
         .Z(n44230)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37335_3_lut.init = 16'hcaca;
    LUT4 i37334_3_lut (.A(\mem[18] [7]), .B(\mem[19] [7]), .C(address[0]), 
         .Z(n44229)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37334_3_lut.init = 16'hcaca;
    LUT4 i37333_3_lut (.A(\mem[16] [7]), .B(\mem[17] [7]), .C(address[0]), 
         .Z(n44228)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37333_3_lut.init = 16'hcaca;
    PFUMX i37657 (.BLUT(n44542), .ALUT(n44543), .C0(address[1]), .Z(n44552));
    LUT4 i37332_3_lut (.A(\mem[14] [7]), .B(\mem[15] [7]), .C(address[0]), 
         .Z(n44227)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37332_3_lut.init = 16'hcaca;
    LUT4 i37331_3_lut (.A(\mem[12] [7]), .B(\mem[13] [7]), .C(address[0]), 
         .Z(n44226)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37331_3_lut.init = 16'hcaca;
    LUT4 i37330_3_lut (.A(\mem[10] [7]), .B(\mem[11] [7]), .C(address[0]), 
         .Z(n44225)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37330_3_lut.init = 16'hcaca;
    PFUMX i37658 (.BLUT(n44544), .ALUT(n44545), .C0(address[1]), .Z(n44553));
    LUT4 i37329_3_lut (.A(\mem[8] [7]), .B(\mem[9] [7]), .C(address[0]), 
         .Z(n44224)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37329_3_lut.init = 16'hcaca;
    LUT4 i37328_3_lut (.A(\mem[6] [7]), .B(\mem[7] [7]), .C(address[0]), 
         .Z(n44223)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37328_3_lut.init = 16'hcaca;
    LUT4 i37327_3_lut (.A(\mem[4] [7]), .B(\mem[5] [7]), .C(address[0]), 
         .Z(n44222)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37327_3_lut.init = 16'hcaca;
    LUT4 i37326_3_lut (.A(\mem[2] [7]), .B(\mem[3] [7]), .C(address[0]), 
         .Z(n44221)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37326_3_lut.init = 16'hcaca;
    LUT4 i37325_3_lut (.A(\mem[0] [7]), .B(\mem[1] [7]), .C(address[0]), 
         .Z(n44220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37325_3_lut.init = 16'hcaca;
    LUT4 i37774_3_lut (.A(\mem[62] [6]), .B(\mem[63] [6]), .C(address[0]), 
         .Z(n44669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37774_3_lut.init = 16'hcaca;
    LUT4 i37773_3_lut (.A(\mem[60] [6]), .B(\mem[61] [6]), .C(address[0]), 
         .Z(n44668)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37773_3_lut.init = 16'hcaca;
    LUT4 i37555_3_lut (.A(\mem[58] [5]), .B(\mem[59] [5]), .C(address[0]), 
         .Z(n44450)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37555_3_lut.init = 16'hcaca;
    LUT4 i37554_3_lut (.A(\mem[56] [5]), .B(\mem[57] [5]), .C(address[0]), 
         .Z(n44449)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37554_3_lut.init = 16'hcaca;
    PFUMX i37465 (.BLUT(n44344), .ALUT(n44345), .C0(address[1]), .Z(n44360));
    LUT4 i37772_3_lut (.A(\mem[58] [6]), .B(\mem[59] [6]), .C(address[0]), 
         .Z(n44667)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37772_3_lut.init = 16'hcaca;
    LUT4 i37771_3_lut (.A(\mem[56] [6]), .B(\mem[57] [6]), .C(address[0]), 
         .Z(n44666)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37771_3_lut.init = 16'hcaca;
    LUT4 i37770_3_lut (.A(\mem[54] [6]), .B(\mem[55] [6]), .C(address[0]), 
         .Z(n44665)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37770_3_lut.init = 16'hcaca;
    PFUMX i37717 (.BLUT(n44600), .ALUT(n44601), .C0(address[1]), .Z(n44612));
    LUT4 i37769_3_lut (.A(\mem[52] [6]), .B(\mem[53] [6]), .C(address[0]), 
         .Z(n44664)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37769_3_lut.init = 16'hcaca;
    LUT4 i37768_3_lut (.A(\mem[50] [6]), .B(\mem[51] [6]), .C(address[0]), 
         .Z(n44663)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37768_3_lut.init = 16'hcaca;
    LUT4 i37767_3_lut (.A(\mem[48] [6]), .B(\mem[49] [6]), .C(address[0]), 
         .Z(n44662)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37767_3_lut.init = 16'hcaca;
    LUT4 i37766_3_lut (.A(\mem[46] [6]), .B(\mem[47] [6]), .C(address[0]), 
         .Z(n44661)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37766_3_lut.init = 16'hcaca;
    LUT4 i37765_3_lut (.A(\mem[44] [6]), .B(\mem[45] [6]), .C(address[0]), 
         .Z(n44660)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37765_3_lut.init = 16'hcaca;
    LUT4 i37764_3_lut (.A(\mem[42] [6]), .B(\mem[43] [6]), .C(address[0]), 
         .Z(n44659)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37764_3_lut.init = 16'hcaca;
    LUT4 i37763_3_lut (.A(\mem[40] [6]), .B(\mem[41] [6]), .C(address[0]), 
         .Z(n44658)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37763_3_lut.init = 16'hcaca;
    LUT4 i37762_3_lut (.A(\mem[38] [6]), .B(\mem[39] [6]), .C(address[0]), 
         .Z(n44657)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37762_3_lut.init = 16'hcaca;
    LUT4 i37761_3_lut (.A(\mem[36] [6]), .B(\mem[37] [6]), .C(address[0]), 
         .Z(n44656)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37761_3_lut.init = 16'hcaca;
    LUT4 i37760_3_lut (.A(\mem[34] [6]), .B(\mem[35] [6]), .C(address[0]), 
         .Z(n44655)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37760_3_lut.init = 16'hcaca;
    LUT4 i37759_3_lut (.A(\mem[32] [6]), .B(\mem[33] [6]), .C(address[0]), 
         .Z(n44654)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37759_3_lut.init = 16'hcaca;
    PFUMX i37466 (.BLUT(n44346), .ALUT(n44347), .C0(address[1]), .Z(n44361));
    LUT4 i37743_3_lut (.A(\mem[62] [7]), .B(\mem[63] [7]), .C(address[0]), 
         .Z(n44638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37743_3_lut.init = 16'hcaca;
    LUT4 i37742_3_lut (.A(\mem[60] [7]), .B(\mem[61] [7]), .C(address[0]), 
         .Z(n44637)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37742_3_lut.init = 16'hcaca;
    LUT4 i37741_3_lut (.A(\mem[58] [7]), .B(\mem[59] [7]), .C(address[0]), 
         .Z(n44636)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37741_3_lut.init = 16'hcaca;
    PFUMX i37467 (.BLUT(n44348), .ALUT(n44349), .C0(address[1]), .Z(n44362));
    LUT4 i37740_3_lut (.A(\mem[56] [7]), .B(\mem[57] [7]), .C(address[0]), 
         .Z(n44635)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37740_3_lut.init = 16'hcaca;
    LUT4 i37739_3_lut (.A(\mem[54] [7]), .B(\mem[55] [7]), .C(address[0]), 
         .Z(n44634)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37739_3_lut.init = 16'hcaca;
    LUT4 i37738_3_lut (.A(\mem[52] [7]), .B(\mem[53] [7]), .C(address[0]), 
         .Z(n44633)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37738_3_lut.init = 16'hcaca;
    LUT4 i37737_3_lut (.A(\mem[50] [7]), .B(\mem[51] [7]), .C(address[0]), 
         .Z(n44632)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37737_3_lut.init = 16'hcaca;
    LUT4 i37736_3_lut (.A(\mem[48] [7]), .B(\mem[49] [7]), .C(address[0]), 
         .Z(n44631)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37736_3_lut.init = 16'hcaca;
    LUT4 i37735_3_lut (.A(\mem[46] [7]), .B(\mem[47] [7]), .C(address[0]), 
         .Z(n44630)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37735_3_lut.init = 16'hcaca;
    LUT4 i37734_3_lut (.A(\mem[44] [7]), .B(\mem[45] [7]), .C(address[0]), 
         .Z(n44629)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37734_3_lut.init = 16'hcaca;
    LUT4 i37733_3_lut (.A(\mem[42] [7]), .B(\mem[43] [7]), .C(address[0]), 
         .Z(n44628)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37733_3_lut.init = 16'hcaca;
    PFUMX i37468 (.BLUT(n44350), .ALUT(n44351), .C0(address[1]), .Z(n44363));
    PFUMX i37469 (.BLUT(n44352), .ALUT(n44353), .C0(address[1]), .Z(n44364));
    LUT4 i37732_3_lut (.A(\mem[40] [7]), .B(\mem[41] [7]), .C(address[0]), 
         .Z(n44627)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37732_3_lut.init = 16'hcaca;
    PFUMX i37470 (.BLUT(n44354), .ALUT(n44355), .C0(address[1]), .Z(n44365));
    LUT4 i37309_3_lut (.A(\mem[30] [6]), .B(\mem[31] [6]), .C(address[0]), 
         .Z(n44204)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37309_3_lut.init = 16'hcaca;
    PFUMX i37471 (.BLUT(n44356), .ALUT(n44357), .C0(address[1]), .Z(n44366));
    LUT4 i37308_3_lut (.A(\mem[28] [6]), .B(\mem[29] [6]), .C(address[0]), 
         .Z(n44203)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37308_3_lut.init = 16'hcaca;
    LUT4 i37731_3_lut (.A(\mem[38] [7]), .B(\mem[39] [7]), .C(address[0]), 
         .Z(n44626)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37731_3_lut.init = 16'hcaca;
    PFUMX i37472 (.BLUT(n44358), .ALUT(n44359), .C0(address[1]), .Z(n44367));
    LUT4 i37730_3_lut (.A(\mem[36] [7]), .B(\mem[37] [7]), .C(address[0]), 
         .Z(n44625)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37730_3_lut.init = 16'hcaca;
    PFUMX i37496 (.BLUT(n44375), .ALUT(n44376), .C0(address[1]), .Z(n44391));
    LUT4 i37307_3_lut (.A(\mem[26] [6]), .B(\mem[27] [6]), .C(address[0]), 
         .Z(n44202)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37307_3_lut.init = 16'hcaca;
    LUT4 i37306_3_lut (.A(\mem[24] [6]), .B(\mem[25] [6]), .C(address[0]), 
         .Z(n44201)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37306_3_lut.init = 16'hcaca;
    PFUMX i37497 (.BLUT(n44377), .ALUT(n44378), .C0(address[1]), .Z(n44392));
    PFUMX i37498 (.BLUT(n44379), .ALUT(n44380), .C0(address[1]), .Z(n44393));
    LUT4 i37729_3_lut (.A(\mem[34] [7]), .B(\mem[35] [7]), .C(address[0]), 
         .Z(n44624)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37729_3_lut.init = 16'hcaca;
    LUT4 i37728_3_lut (.A(\mem[32] [7]), .B(\mem[33] [7]), .C(address[0]), 
         .Z(n44623)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37728_3_lut.init = 16'hcaca;
    LUT4 i37305_3_lut (.A(\mem[22] [6]), .B(\mem[23] [6]), .C(address[0]), 
         .Z(n44200)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37305_3_lut.init = 16'hcaca;
    LUT4 i37304_3_lut (.A(\mem[20] [6]), .B(\mem[21] [6]), .C(address[0]), 
         .Z(n44199)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37304_3_lut.init = 16'hcaca;
    LUT4 i37303_3_lut (.A(\mem[18] [6]), .B(\mem[19] [6]), .C(address[0]), 
         .Z(n44198)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37303_3_lut.init = 16'hcaca;
    LUT4 i37302_3_lut (.A(\mem[16] [6]), .B(\mem[17] [6]), .C(address[0]), 
         .Z(n44197)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37302_3_lut.init = 16'hcaca;
    PFUMX i37499 (.BLUT(n44381), .ALUT(n44382), .C0(address[1]), .Z(n44394));
    LUT4 i37301_3_lut (.A(\mem[14] [6]), .B(\mem[15] [6]), .C(address[0]), 
         .Z(n44196)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37301_3_lut.init = 16'hcaca;
    LUT4 i37300_3_lut (.A(\mem[12] [6]), .B(\mem[13] [6]), .C(address[0]), 
         .Z(n44195)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37300_3_lut.init = 16'hcaca;
    LUT4 i37299_3_lut (.A(\mem[10] [6]), .B(\mem[11] [6]), .C(address[0]), 
         .Z(n44194)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37299_3_lut.init = 16'hcaca;
    LUT4 i37298_3_lut (.A(\mem[8] [6]), .B(\mem[9] [6]), .C(address[0]), 
         .Z(n44193)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37298_3_lut.init = 16'hcaca;
    PFUMX i37500 (.BLUT(n44383), .ALUT(n44384), .C0(address[1]), .Z(n44395));
    LUT4 i37297_3_lut (.A(\mem[6] [6]), .B(\mem[7] [6]), .C(address[0]), 
         .Z(n44192)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37297_3_lut.init = 16'hcaca;
    PFUMX i37501 (.BLUT(n44385), .ALUT(n44386), .C0(address[1]), .Z(n44396));
    PFUMX i37502 (.BLUT(n44387), .ALUT(n44388), .C0(address[1]), .Z(n44397));
    LUT4 i37296_3_lut (.A(\mem[4] [6]), .B(\mem[5] [6]), .C(address[0]), 
         .Z(n44191)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37296_3_lut.init = 16'hcaca;
    PFUMX i37503 (.BLUT(n44389), .ALUT(n44390), .C0(address[1]), .Z(n44398));
    PFUMX i37682 (.BLUT(n44561), .ALUT(n44562), .C0(address[1]), .Z(n44577));
    LUT4 i37295_3_lut (.A(\mem[2] [6]), .B(\mem[3] [6]), .C(address[0]), 
         .Z(n44190)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37295_3_lut.init = 16'hcaca;
    LUT4 i37294_3_lut (.A(\mem[0] [6]), .B(\mem[1] [6]), .C(address[0]), 
         .Z(n44189)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37294_3_lut.init = 16'hcaca;
    PFUMX i37683 (.BLUT(n44563), .ALUT(n44564), .C0(address[1]), .Z(n44578));
    PFUMX i37684 (.BLUT(n44565), .ALUT(n44566), .C0(address[1]), .Z(n44579));
    PFUMX i37685 (.BLUT(n44567), .ALUT(n44568), .C0(address[1]), .Z(n44580));
    LUT4 i37553_3_lut (.A(\mem[54] [5]), .B(\mem[55] [5]), .C(address[0]), 
         .Z(n44448)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37553_3_lut.init = 16'hcaca;
    PFUMX i37686 (.BLUT(n44569), .ALUT(n44570), .C0(address[1]), .Z(n44581));
    PFUMX i37687 (.BLUT(n44571), .ALUT(n44572), .C0(address[1]), .Z(n44582));
    PFUMX i37688 (.BLUT(n44573), .ALUT(n44574), .C0(address[1]), .Z(n44583));
    LUT4 i37552_3_lut (.A(\mem[52] [5]), .B(\mem[53] [5]), .C(address[0]), 
         .Z(n44447)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37552_3_lut.init = 16'hcaca;
    PFUMX i37527 (.BLUT(n44406), .ALUT(n44407), .C0(address[1]), .Z(n44422));
    PFUMX i37528 (.BLUT(n44408), .ALUT(n44409), .C0(address[1]), .Z(n44423));
    PFUMX i37529 (.BLUT(n44410), .ALUT(n44411), .C0(address[1]), .Z(n44424));
    PFUMX i37689 (.BLUT(n44575), .ALUT(n44576), .C0(address[1]), .Z(n44584));
    PFUMX i37530 (.BLUT(n44412), .ALUT(n44413), .C0(address[1]), .Z(n44425));
    LUT4 Select_6139_i3_3_lut_4_lut (.A(akku_o_c_4), .B(n46211), .C(data_7__N_102), 
         .D(data_7__N_89[4]), .Z(data[4])) /* synthesis lut_function=(A ((C (D))+!B)+!A (C (D))) */ ;
    defparam Select_6139_i3_3_lut_4_lut.init = 16'hf222;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n46211), .B(n46856), .C(n43653), .D(n46220), 
         .Z(mem_62__7__N_294)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_8 (.A(n46211), .B(n46856), .C(n46239), 
         .D(n46237), .Z(mem_39__7__N_225)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_8.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_9 (.A(n46211), .B(n46856), .C(n46238), 
         .D(n46237), .Z(mem_31__7__N_201)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_9.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_10 (.A(n46211), .B(n46856), .C(n43635), 
         .D(n46242), .Z(mem_53__7__N_267)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_10.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_11 (.A(n46211), .B(n46856), .C(n43636), 
         .D(n46242), .Z(mem_52__7__N_264)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_11.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_12 (.A(n46211), .B(n46856), .C(n23757), 
         .D(n46242), .Z(mem_51__7__N_261)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_12.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_13 (.A(n46211), .B(n46856), .C(n43654), 
         .D(n46242), .Z(mem_50__7__N_258)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_13.init = 16'h0004;
    LUT4 i2_3_lut_rep_1051_4_lut (.A(n46211), .B(n46856), .C(address[2]), 
         .D(address[1]), .Z(n46172)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i2_3_lut_rep_1051_4_lut.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_14 (.A(n46211), .B(n46856), .C(n46220), 
         .D(n46237), .Z(mem_63__7__N_297)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_14.init = 16'h4000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_15 (.A(n46211), .B(n46856), .C(n46242), 
         .D(n46237), .Z(mem_55__7__N_273)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_15.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_16 (.A(n46211), .B(n46856), .C(n46241), 
         .D(n46237), .Z(mem_47__7__N_249)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_16.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_17 (.A(n46211), .B(n46856), .C(n46234), 
         .D(n46237), .Z(mem_15__7__N_153)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_17.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_18 (.A(n46211), .B(n46856), .C(n43653), 
         .D(n46242), .Z(mem_54__7__N_270)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_18.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_19 (.A(n46211), .B(n46856), .C(n43654), 
         .D(n46241), .Z(mem_42__7__N_234)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_19.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_20 (.A(n46211), .B(n46856), .C(n23757), 
         .D(n46241), .Z(mem_43__7__N_237)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_20.init = 16'h0004;
    PFUMX i37531 (.BLUT(n44414), .ALUT(n44415), .C0(address[1]), .Z(n44426));
    LUT4 i1_2_lut_3_lut_4_lut_adj_21 (.A(n46211), .B(n46856), .C(n43636), 
         .D(n46241), .Z(mem_44__7__N_240)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_21.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_22 (.A(n46211), .B(n46856), .C(n43635), 
         .D(n46241), .Z(mem_45__7__N_243)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_22.init = 16'h0004;
    PFUMX i37532 (.BLUT(n44416), .ALUT(n44417), .C0(address[1]), .Z(n44427));
    LUT4 i1_2_lut_3_lut_4_lut_adj_23 (.A(n46211), .B(n46856), .C(n43653), 
         .D(n46241), .Z(mem_46__7__N_246)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_23.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_24 (.A(n46211), .B(n46856), .C(n43654), 
         .D(n46239), .Z(mem_34__7__N_210)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_24.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_25 (.A(n46211), .B(n46856), .C(n23757), 
         .D(n46239), .Z(mem_35__7__N_213)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_25.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_26 (.A(n46211), .B(n46856), .C(n43636), 
         .D(n46239), .Z(mem_36__7__N_216)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_26.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_27 (.A(n46211), .B(n46856), .C(n43635), 
         .D(n46239), .Z(mem_37__7__N_219)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_27.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_28 (.A(n46211), .B(n46856), .C(n43653), 
         .D(n46239), .Z(mem_38__7__N_222)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_28.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_29 (.A(n46211), .B(n46856), .C(n43654), 
         .D(n46238), .Z(mem_26__7__N_186)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_29.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_30 (.A(n46211), .B(n46856), .C(n23757), 
         .D(n46238), .Z(mem_27__7__N_189)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_30.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_31 (.A(n46211), .B(n46856), .C(n43636), 
         .D(n46238), .Z(mem_28__7__N_192)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_31.init = 16'h0004;
    PFUMX i37533 (.BLUT(n44418), .ALUT(n44419), .C0(address[1]), .Z(n44428));
    LUT4 i1_2_lut_3_lut_4_lut_adj_32 (.A(n46211), .B(n46856), .C(n43635), 
         .D(n46238), .Z(mem_29__7__N_195)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_32.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_33 (.A(n46211), .B(n46856), .C(n43653), 
         .D(n46238), .Z(mem_30__7__N_198)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_33.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_34 (.A(n46211), .B(n46856), .C(n43654), 
         .D(n46236), .Z(mem_18__7__N_162)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_34.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_35 (.A(n46211), .B(n46856), .C(n23757), 
         .D(n46236), .Z(mem_19__7__N_165)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_35.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_36 (.A(n46211), .B(n46856), .C(n43636), 
         .D(n46236), .Z(mem_20__7__N_168)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_36.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_37 (.A(n46211), .B(n46856), .C(n43635), 
         .D(n46236), .Z(mem_21__7__N_171)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_37.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_38 (.A(n46211), .B(n46856), .C(n43653), 
         .D(n46236), .Z(mem_22__7__N_174)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_38.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_39 (.A(n46211), .B(n46856), .C(n46237), 
         .D(n46236), .Z(mem_23__7__N_177)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_39.init = 16'h0040;
    LUT4 i1_2_lut_3_lut_4_lut_adj_40 (.A(n46211), .B(n46856), .C(n43654), 
         .D(n46234), .Z(mem_10__7__N_138)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_40.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_41 (.A(n46211), .B(n46856), .C(n23757), 
         .D(n46234), .Z(mem_11__7__N_141)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_41.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_42 (.A(n46211), .B(n46856), .C(n43636), 
         .D(n46234), .Z(mem_12__7__N_144)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_42.init = 16'h0004;
    PFUMX i37534 (.BLUT(n44420), .ALUT(n44421), .C0(address[1]), .Z(n44429));
    LUT4 i1_2_lut_3_lut_4_lut_adj_43 (.A(n46211), .B(n46856), .C(n43635), 
         .D(n46234), .Z(mem_13__7__N_147)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_43.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_44 (.A(n46211), .B(n46856), .C(n43653), 
         .D(n46234), .Z(mem_14__7__N_150)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_44.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_45 (.A(n46211), .B(n46856), .C(n43635), 
         .D(n46220), .Z(mem_61__7__N_291)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_45.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_46 (.A(n46211), .B(n46856), .C(n43636), 
         .D(n46220), .Z(mem_60__7__N_288)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_46.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_47 (.A(n46211), .B(n46856), .C(n43654), 
         .D(n46232), .Z(mem_2__7__N_114)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_47.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_48 (.A(n46211), .B(n46856), .C(n23757), 
         .D(n46220), .Z(mem_59__7__N_285)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_48.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_49 (.A(n46211), .B(n46856), .C(n43654), 
         .D(n46220), .Z(mem_58__7__N_282)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_49.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_50 (.A(n46211), .B(n46856), .C(n46237), 
         .D(n46232), .Z(mem_7__7__N_129)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_50.init = 16'h0040;
    LUT4 i1_2_lut_3_lut_4_lut_adj_51 (.A(n46211), .B(n46856), .C(n43653), 
         .D(n46232), .Z(mem_6__7__N_126)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_51.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_52 (.A(n46211), .B(n46856), .C(n43635), 
         .D(n46232), .Z(mem_5__7__N_123)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_52.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_53 (.A(n46211), .B(n46856), .C(n43636), 
         .D(n46232), .Z(mem_4__7__N_120)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_53.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut_adj_54 (.A(n46211), .B(n46856), .C(n23757), 
         .D(n46232), .Z(mem_3__7__N_117)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_3_lut_4_lut_adj_54.init = 16'h0004;
    LUT4 Select_6143_i3_3_lut_4_lut (.A(akku_o_c_0), .B(n46211), .C(data_7__N_102), 
         .D(data_7__N_89[0]), .Z(data[0])) /* synthesis lut_function=(A ((C (D))+!B)+!A (C (D))) */ ;
    defparam Select_6143_i3_3_lut_4_lut.init = 16'hf222;
    PFUMX i37718 (.BLUT(n44602), .ALUT(n44603), .C0(address[1]), .Z(n44613));
    LUT4 i37789_3_lut (.A(n44682), .B(n44683), .C(address[4]), .Z(n44684)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37789_3_lut.init = 16'hcaca;
    LUT4 i37324_3_lut (.A(n44217), .B(n44218), .C(address[4]), .Z(n44219)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37324_3_lut.init = 16'hcaca;
    LUT4 i37758_3_lut (.A(n44651), .B(n44652), .C(address[4]), .Z(n44653)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37758_3_lut.init = 16'hcaca;
    LUT4 i37355_3_lut (.A(n44248), .B(n44249), .C(address[4]), .Z(n44250)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37355_3_lut.init = 16'hcaca;
    LUT4 i37727_3_lut (.A(n44620), .B(n44621), .C(address[4]), .Z(n44622)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37727_3_lut.init = 16'hcaca;
    LUT4 i37386_3_lut (.A(n44279), .B(n44280), .C(address[4]), .Z(n44281)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37386_3_lut.init = 16'hcaca;
    LUT4 i37696_3_lut (.A(n44589), .B(n44590), .C(address[4]), .Z(n44591)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37696_3_lut.init = 16'hcaca;
    LUT4 i37417_3_lut (.A(n44310), .B(n44311), .C(address[4]), .Z(n44312)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37417_3_lut.init = 16'hcaca;
    LUT4 Select_6136_i3_3_lut_4_lut (.A(akku_o_c_7), .B(n46211), .C(data_7__N_102), 
         .D(data_7__N_89[7]), .Z(data[7])) /* synthesis lut_function=(A ((C (D))+!B)+!A (C (D))) */ ;
    defparam Select_6136_i3_3_lut_4_lut.init = 16'hf222;
    LUT4 Select_6137_i3_3_lut_4_lut (.A(akku_o_c_6), .B(n46211), .C(data_7__N_102), 
         .D(data_7__N_89[6]), .Z(data[6])) /* synthesis lut_function=(A ((C (D))+!B)+!A (C (D))) */ ;
    defparam Select_6137_i3_3_lut_4_lut.init = 16'hf222;
    PFUMX i37558 (.BLUT(n44437), .ALUT(n44438), .C0(address[1]), .Z(n44453));
    LUT4 i37665_3_lut (.A(n44558), .B(n44559), .C(address[4]), .Z(n44560)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37665_3_lut.init = 16'hcaca;
    PFUMX i37719 (.BLUT(n44604), .ALUT(n44605), .C0(address[1]), .Z(n44614));
    LUT4 Select_6138_i3_3_lut_4_lut (.A(akku_o_c_5), .B(n46211), .C(data_7__N_102), 
         .D(data_7__N_89[5]), .Z(data[5])) /* synthesis lut_function=(A ((C (D))+!B)+!A (C (D))) */ ;
    defparam Select_6138_i3_3_lut_4_lut.init = 16'hf222;
    LUT4 Select_6140_i3_3_lut_4_lut (.A(akku_o_c_3), .B(n46211), .C(data_7__N_102), 
         .D(data_7__N_89[3]), .Z(data[3])) /* synthesis lut_function=(A ((C (D))+!B)+!A (C (D))) */ ;
    defparam Select_6140_i3_3_lut_4_lut.init = 16'hf222;
    LUT4 Select_6141_i3_3_lut_4_lut (.A(akku_o_c_2), .B(n46211), .C(data_7__N_102), 
         .D(data_7__N_89[2]), .Z(data[2])) /* synthesis lut_function=(A ((C (D))+!B)+!A (C (D))) */ ;
    defparam Select_6141_i3_3_lut_4_lut.init = 16'hf222;
    LUT4 Select_6142_i3_3_lut_4_lut (.A(akku_o_c_1), .B(n46211), .C(data_7__N_102), 
         .D(data_7__N_89[1]), .Z(data[1])) /* synthesis lut_function=(A ((C (D))+!B)+!A (C (D))) */ ;
    defparam Select_6142_i3_3_lut_4_lut.init = 16'hf222;
    LUT4 i37448_3_lut (.A(n44341), .B(n44342), .C(address[4]), .Z(n44343)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37448_3_lut.init = 16'hcaca;
    LUT4 i37634_3_lut (.A(n44527), .B(n44528), .C(address[4]), .Z(n44529)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37634_3_lut.init = 16'hcaca;
    LUT4 i37479_3_lut (.A(n44372), .B(n44373), .C(address[4]), .Z(n44374)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37479_3_lut.init = 16'hcaca;
    LUT4 i37603_3_lut (.A(n44496), .B(n44497), .C(address[4]), .Z(n44498)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37603_3_lut.init = 16'hcaca;
    LUT4 i37510_3_lut (.A(n44403), .B(n44404), .C(address[4]), .Z(n44405)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37510_3_lut.init = 16'hcaca;
    LUT4 i37572_3_lut (.A(n44465), .B(n44466), .C(address[4]), .Z(n44467)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37572_3_lut.init = 16'hcaca;
    LUT4 i37541_3_lut (.A(n44434), .B(n44435), .C(address[4]), .Z(n44436)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37541_3_lut.init = 16'hcaca;
    PFUMX i37559 (.BLUT(n44439), .ALUT(n44440), .C0(address[1]), .Z(n44454));
    PFUMX i37560 (.BLUT(n44441), .ALUT(n44442), .C0(address[1]), .Z(n44455));
    PFUMX i37561 (.BLUT(n44443), .ALUT(n44444), .C0(address[1]), .Z(n44456));
    LUT4 i1_2_lut_3_lut_4_lut_adj_55 (.A(address[3]), .B(n46278), .C(address[0]), 
         .D(n46172), .Z(mem_57__7__N_279)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_55.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_56 (.A(address[3]), .B(n46278), .C(address[0]), 
         .D(n46172), .Z(mem_56__7__N_276)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_56.init = 16'h0800;
    LUT4 i37551_3_lut (.A(\mem[50] [5]), .B(\mem[51] [5]), .C(address[0]), 
         .Z(n44446)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37551_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_57 (.A(address[5]), .B(n46274), .C(address[0]), 
         .D(n46172), .Z(mem_0__7__N_106)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_57.init = 16'h0100;
    LUT4 i1_2_lut_3_lut_4_lut_adj_58 (.A(address[5]), .B(n46274), .C(address[0]), 
         .D(n46172), .Z(mem_1__7__N_111)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_58.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_59 (.A(address[5]), .B(n46275), .C(address[0]), 
         .D(n46172), .Z(mem_8__7__N_132)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_59.init = 16'h0100;
    LUT4 i1_2_lut_3_lut_4_lut_adj_60 (.A(address[5]), .B(n46275), .C(address[0]), 
         .D(n46172), .Z(mem_9__7__N_135)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_60.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_61 (.A(address[3]), .B(n46273), .C(address[0]), 
         .D(n46172), .Z(mem_16__7__N_156)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_61.init = 16'h0100;
    LUT4 i1_2_lut_3_lut_4_lut_adj_62 (.A(address[3]), .B(n46273), .C(address[0]), 
         .D(n46172), .Z(mem_17__7__N_159)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_62.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_63 (.A(address[3]), .B(n46273), .C(address[0]), 
         .D(n46172), .Z(mem_24__7__N_180)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_63.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_64 (.A(address[3]), .B(n46273), .C(address[0]), 
         .D(n46172), .Z(mem_25__7__N_183)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_64.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_65 (.A(address[5]), .B(n46274), .C(address[0]), 
         .D(n46172), .Z(mem_32__7__N_204)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_65.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_66 (.A(address[5]), .B(n46274), .C(address[0]), 
         .D(n46172), .Z(mem_33__7__N_207)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_66.init = 16'h2000;
    PFUMX i37720 (.BLUT(n44606), .ALUT(n44607), .C0(address[1]), .Z(n44615));
    LUT4 i1_2_lut_3_lut_4_lut_adj_67 (.A(address[5]), .B(n46275), .C(address[0]), 
         .D(n46172), .Z(mem_40__7__N_228)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_67.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_68 (.A(address[5]), .B(n46275), .C(address[0]), 
         .D(n46172), .Z(mem_41__7__N_231)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_68.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_69 (.A(address[3]), .B(n46278), .C(address[0]), 
         .D(n46172), .Z(mem_48__7__N_252)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_69.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_70 (.A(address[3]), .B(n46278), .C(address[0]), 
         .D(n46172), .Z(mem_49__7__N_255)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_4_lut_adj_70.init = 16'h4000;
    LUT4 i1_2_lut_rep_1170 (.A(reset_c), .B(clk_c), .Z(n46856)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_2_lut_rep_1170.init = 16'h2222;
    LUT4 i1_4_lut_4_lut_4_lut_3_lut_4_lut (.A(reset_c), .B(clk_c), .C(\states[0] ), 
         .D(\states[1] ), .Z(data_7__N_102)) /* synthesis lut_function=(!((B+!((D)+!C))+!A)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(65[13] 78[20])
    defparam i1_4_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h2202;
    LUT4 i1_2_lut_3_lut (.A(address[0]), .B(address[1]), .C(address[2]), 
         .Z(n43653)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut.init = 16'hbfbf;
    LUT4 i1_2_lut_3_lut_adj_71 (.A(address[0]), .B(address[1]), .C(address[2]), 
         .Z(n43654)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_adj_71.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_adj_72 (.A(address[1]), .B(address[2]), .C(address[0]), 
         .Z(n43635)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_adj_72.init = 16'hbfbf;
    LUT4 i1_2_lut_3_lut_adj_73 (.A(address[1]), .B(address[2]), .C(address[0]), 
         .Z(n43636)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/10352/vhdl-labs/lab9_mcpu/sram64kx8.vhd(67[22:29])
    defparam i1_2_lut_3_lut_adj_73.init = 16'hfbfb;
    LUT4 i23741_2_lut_rep_1157 (.A(address[4]), .B(address[5]), .Z(n46278)) /* synthesis lut_function=(A (B)) */ ;
    defparam i23741_2_lut_rep_1157.init = 16'h8888;
    LUT4 i24261_2_lut_rep_1099_3_lut (.A(address[4]), .B(address[5]), .C(address[3]), 
         .Z(n46220)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i24261_2_lut_rep_1099_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_1121_3_lut (.A(address[4]), .B(address[5]), .C(address[3]), 
         .Z(n46242)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_rep_1121_3_lut.init = 16'hf7f7;
    LUT4 i37550_3_lut (.A(\mem[48] [5]), .B(\mem[49] [5]), .C(address[0]), 
         .Z(n44445)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37550_3_lut.init = 16'hcaca;
    
endmodule
